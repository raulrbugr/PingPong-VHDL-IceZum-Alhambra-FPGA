// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Mar 17 2018 18:15:53

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "incremental" view "INTERFACE"

module incremental (
    leds,
    reset,
    clk);

    output [7:0] leds;
    input reset;
    input clk;

    wire N__2704;
    wire N__2703;
    wire N__2702;
    wire N__2694;
    wire N__2693;
    wire N__2692;
    wire N__2683;
    wire N__2682;
    wire N__2681;
    wire N__2674;
    wire N__2673;
    wire N__2672;
    wire N__2665;
    wire N__2664;
    wire N__2663;
    wire N__2656;
    wire N__2655;
    wire N__2654;
    wire N__2647;
    wire N__2646;
    wire N__2645;
    wire N__2638;
    wire N__2637;
    wire N__2636;
    wire N__2629;
    wire N__2628;
    wire N__2627;
    wire N__2620;
    wire N__2619;
    wire N__2618;
    wire N__2601;
    wire N__2598;
    wire N__2595;
    wire N__2594;
    wire N__2591;
    wire N__2588;
    wire N__2587;
    wire N__2584;
    wire N__2579;
    wire N__2574;
    wire N__2571;
    wire N__2570;
    wire N__2567;
    wire N__2564;
    wire N__2563;
    wire N__2560;
    wire N__2555;
    wire N__2550;
    wire N__2547;
    wire N__2544;
    wire N__2541;
    wire N__2540;
    wire N__2539;
    wire N__2536;
    wire N__2531;
    wire N__2526;
    wire N__2525;
    wire N__2524;
    wire N__2523;
    wire N__2522;
    wire N__2521;
    wire N__2520;
    wire N__2505;
    wire N__2504;
    wire N__2503;
    wire N__2502;
    wire N__2501;
    wire N__2498;
    wire N__2491;
    wire N__2490;
    wire N__2487;
    wire N__2484;
    wire N__2481;
    wire N__2478;
    wire N__2469;
    wire N__2468;
    wire N__2467;
    wire N__2462;
    wire N__2459;
    wire N__2454;
    wire N__2451;
    wire N__2448;
    wire N__2447;
    wire N__2446;
    wire N__2443;
    wire N__2438;
    wire N__2433;
    wire N__2430;
    wire N__2427;
    wire N__2424;
    wire N__2423;
    wire N__2420;
    wire N__2417;
    wire N__2416;
    wire N__2413;
    wire N__2408;
    wire N__2403;
    wire N__2400;
    wire N__2397;
    wire N__2396;
    wire N__2393;
    wire N__2390;
    wire N__2387;
    wire N__2384;
    wire N__2379;
    wire N__2378;
    wire N__2377;
    wire N__2376;
    wire N__2373;
    wire N__2372;
    wire N__2371;
    wire N__2370;
    wire N__2363;
    wire N__2354;
    wire N__2351;
    wire N__2350;
    wire N__2349;
    wire N__2348;
    wire N__2347;
    wire N__2346;
    wire N__2345;
    wire N__2344;
    wire N__2343;
    wire N__2342;
    wire N__2341;
    wire N__2340;
    wire N__2339;
    wire N__2338;
    wire N__2337;
    wire N__2336;
    wire N__2333;
    wire N__2330;
    wire N__2321;
    wire N__2312;
    wire N__2305;
    wire N__2296;
    wire N__2283;
    wire N__2280;
    wire N__2277;
    wire N__2276;
    wire N__2275;
    wire N__2272;
    wire N__2269;
    wire N__2266;
    wire N__2263;
    wire N__2260;
    wire N__2253;
    wire N__2252;
    wire N__2247;
    wire N__2246;
    wire N__2245;
    wire N__2244;
    wire N__2243;
    wire N__2242;
    wire N__2241;
    wire N__2240;
    wire N__2239;
    wire N__2238;
    wire N__2237;
    wire N__2236;
    wire N__2235;
    wire N__2234;
    wire N__2233;
    wire N__2230;
    wire N__2215;
    wire N__2214;
    wire N__2199;
    wire N__2198;
    wire N__2197;
    wire N__2196;
    wire N__2195;
    wire N__2194;
    wire N__2193;
    wire N__2192;
    wire N__2189;
    wire N__2186;
    wire N__2183;
    wire N__2180;
    wire N__2175;
    wire N__2164;
    wire N__2151;
    wire N__2148;
    wire N__2145;
    wire N__2142;
    wire N__2141;
    wire N__2140;
    wire N__2137;
    wire N__2134;
    wire N__2131;
    wire N__2128;
    wire N__2125;
    wire N__2118;
    wire N__2117;
    wire N__2116;
    wire N__2115;
    wire N__2114;
    wire N__2113;
    wire N__2112;
    wire N__2111;
    wire N__2110;
    wire N__2091;
    wire N__2088;
    wire N__2085;
    wire N__2084;
    wire N__2083;
    wire N__2082;
    wire N__2081;
    wire N__2070;
    wire N__2067;
    wire N__2064;
    wire N__2063;
    wire N__2062;
    wire N__2061;
    wire N__2060;
    wire N__2059;
    wire N__2058;
    wire N__2057;
    wire N__2056;
    wire N__2037;
    wire N__2034;
    wire N__2031;
    wire N__2030;
    wire N__2027;
    wire N__2026;
    wire N__2023;
    wire N__2020;
    wire N__2017;
    wire N__2010;
    wire N__2007;
    wire N__2004;
    wire N__2001;
    wire N__2000;
    wire N__1999;
    wire N__1996;
    wire N__1993;
    wire N__1990;
    wire N__1983;
    wire N__1980;
    wire N__1977;
    wire N__1974;
    wire N__1971;
    wire N__1970;
    wire N__1967;
    wire N__1964;
    wire N__1961;
    wire N__1956;
    wire N__1953;
    wire N__1950;
    wire N__1947;
    wire N__1946;
    wire N__1945;
    wire N__1942;
    wire N__1937;
    wire N__1932;
    wire N__1929;
    wire N__1928;
    wire N__1927;
    wire N__1922;
    wire N__1919;
    wire N__1914;
    wire N__1911;
    wire N__1908;
    wire N__1907;
    wire N__1906;
    wire N__1903;
    wire N__1900;
    wire N__1897;
    wire N__1890;
    wire N__1887;
    wire N__1884;
    wire N__1881;
    wire N__1880;
    wire N__1879;
    wire N__1876;
    wire N__1873;
    wire N__1870;
    wire N__1863;
    wire N__1862;
    wire N__1861;
    wire N__1858;
    wire N__1855;
    wire N__1852;
    wire N__1849;
    wire N__1842;
    wire N__1839;
    wire N__1836;
    wire N__1833;
    wire N__1832;
    wire N__1831;
    wire N__1828;
    wire N__1825;
    wire N__1822;
    wire N__1819;
    wire N__1816;
    wire N__1809;
    wire N__1806;
    wire N__1803;
    wire N__1800;
    wire N__1799;
    wire N__1798;
    wire N__1795;
    wire N__1792;
    wire N__1789;
    wire N__1786;
    wire N__1779;
    wire N__1776;
    wire N__1773;
    wire N__1770;
    wire N__1769;
    wire N__1768;
    wire N__1765;
    wire N__1762;
    wire N__1759;
    wire N__1756;
    wire N__1749;
    wire N__1746;
    wire N__1743;
    wire N__1740;
    wire N__1739;
    wire N__1736;
    wire N__1735;
    wire N__1732;
    wire N__1729;
    wire N__1726;
    wire N__1719;
    wire N__1716;
    wire N__1713;
    wire N__1710;
    wire N__1709;
    wire N__1708;
    wire N__1705;
    wire N__1702;
    wire N__1699;
    wire N__1696;
    wire N__1693;
    wire N__1686;
    wire N__1683;
    wire N__1680;
    wire N__1677;
    wire N__1676;
    wire N__1673;
    wire N__1672;
    wire N__1669;
    wire N__1666;
    wire N__1663;
    wire N__1656;
    wire N__1653;
    wire N__1650;
    wire N__1647;
    wire N__1646;
    wire N__1645;
    wire N__1642;
    wire N__1639;
    wire N__1636;
    wire N__1633;
    wire N__1626;
    wire N__1623;
    wire N__1620;
    wire N__1617;
    wire N__1616;
    wire N__1615;
    wire N__1612;
    wire N__1609;
    wire N__1606;
    wire N__1603;
    wire N__1596;
    wire N__1593;
    wire N__1590;
    wire N__1587;
    wire N__1586;
    wire N__1585;
    wire N__1582;
    wire N__1579;
    wire N__1576;
    wire N__1573;
    wire N__1570;
    wire N__1563;
    wire N__1560;
    wire N__1557;
    wire N__1554;
    wire N__1553;
    wire N__1552;
    wire N__1549;
    wire N__1546;
    wire N__1543;
    wire N__1540;
    wire N__1533;
    wire N__1530;
    wire N__1527;
    wire N__1524;
    wire N__1523;
    wire N__1522;
    wire N__1519;
    wire N__1516;
    wire N__1513;
    wire N__1510;
    wire N__1503;
    wire N__1500;
    wire N__1497;
    wire N__1494;
    wire N__1491;
    wire N__1490;
    wire N__1489;
    wire N__1486;
    wire N__1483;
    wire N__1480;
    wire N__1477;
    wire N__1474;
    wire N__1467;
    wire N__1464;
    wire N__1461;
    wire N__1458;
    wire N__1455;
    wire N__1454;
    wire N__1453;
    wire N__1450;
    wire N__1447;
    wire N__1444;
    wire N__1441;
    wire N__1434;
    wire N__1431;
    wire N__1428;
    wire N__1425;
    wire N__1424;
    wire N__1419;
    wire N__1416;
    wire N__1413;
    wire N__1410;
    wire N__1409;
    wire N__1404;
    wire N__1401;
    wire N__1400;
    wire N__1399;
    wire N__1396;
    wire N__1393;
    wire N__1390;
    wire N__1383;
    wire N__1382;
    wire N__1381;
    wire N__1378;
    wire N__1375;
    wire N__1372;
    wire N__1365;
    wire N__1364;
    wire N__1363;
    wire N__1360;
    wire N__1357;
    wire N__1354;
    wire N__1351;
    wire N__1344;
    wire N__1341;
    wire N__1338;
    wire N__1335;
    wire N__1334;
    wire N__1333;
    wire N__1330;
    wire N__1327;
    wire N__1324;
    wire N__1321;
    wire N__1318;
    wire N__1311;
    wire N__1308;
    wire N__1305;
    wire N__1302;
    wire N__1301;
    wire N__1300;
    wire N__1297;
    wire N__1294;
    wire N__1291;
    wire N__1288;
    wire N__1281;
    wire N__1278;
    wire N__1275;
    wire N__1272;
    wire N__1271;
    wire N__1270;
    wire N__1267;
    wire N__1264;
    wire N__1261;
    wire N__1258;
    wire N__1251;
    wire N__1248;
    wire N__1245;
    wire N__1242;
    wire N__1241;
    wire N__1240;
    wire N__1237;
    wire N__1234;
    wire N__1231;
    wire N__1224;
    wire N__1223;
    wire N__1220;
    wire N__1217;
    wire N__1212;
    wire N__1211;
    wire N__1210;
    wire N__1207;
    wire N__1204;
    wire N__1203;
    wire N__1194;
    wire N__1191;
    wire N__1190;
    wire N__1189;
    wire N__1186;
    wire N__1185;
    wire N__1180;
    wire N__1175;
    wire N__1170;
    wire N__1169;
    wire N__1168;
    wire N__1163;
    wire N__1160;
    wire N__1155;
    wire N__1154;
    wire N__1153;
    wire N__1150;
    wire N__1145;
    wire N__1142;
    wire N__1137;
    wire N__1134;
    wire N__1131;
    wire N__1128;
    wire N__1125;
    wire N__1122;
    wire N__1119;
    wire N__1116;
    wire N__1113;
    wire N__1110;
    wire N__1107;
    wire N__1104;
    wire N__1101;
    wire N__1098;
    wire N__1095;
    wire N__1092;
    wire GNDG0;
    wire VCCG0;
    wire op_eq_un4_fin_cnt_20_3_cascade_;
    wire op_eq_un4_fin_cnt_20_4;
    wire op_eq_un4_fin_cnt_21_9;
    wire op_eq_un4_fin_cnt_21_11;
    wire op_eq_un4_fin_cnt_21_10;
    wire op_eq_un4_fin_cnt_21_8;
    wire op_eq_un4_fin_cnt_20;
    wire op_eq_un4_fin_cnt_21;
    wire \UC.epZ0Z_3 ;
    wire \UC.epZ0Z_6 ;
    wire \UC.value_cnte_0_i ;
    wire \UC.epZ0Z_4 ;
    wire \UC.sr_reg ;
    wire \UC.epZ0Z_0 ;
    wire \UC.epZ0Z_8 ;
    wire \UC.epZ0Z_1 ;
    wire \UC.epZ0Z_7 ;
    wire value_cntZ0Z_0;
    wire bfn_6_5_0_;
    wire value_cntZ0Z_1;
    wire value_cnt_cry_0_THRU_CO;
    wire value_cnt_cry_0;
    wire value_cntZ0Z_2;
    wire value_cnt_cry_1_THRU_CO;
    wire value_cnt_cry_1;
    wire value_cntZ0Z_3;
    wire value_cnt_cry_2_THRU_CO;
    wire value_cnt_cry_2;
    wire value_cntZ0Z_4;
    wire value_cnt_cry_3_THRU_CO;
    wire value_cnt_cry_3;
    wire value_cntZ0Z_5;
    wire value_cnt_cry_4_THRU_CO;
    wire value_cnt_cry_4;
    wire value_cntZ0Z_6;
    wire value_cnt_cry_5_THRU_CO;
    wire value_cnt_cry_5;
    wire value_cntZ0Z_7;
    wire value_cnt_cry_6_THRU_CO;
    wire value_cnt_cry_6;
    wire value_cnt_cry_7;
    wire value_cntZ0Z_8;
    wire value_cnt_cry_7_THRU_CO;
    wire bfn_6_6_0_;
    wire value_cnt_cry_8;
    wire value_cntZ0Z_10;
    wire value_cnt_cry_9_THRU_CO;
    wire value_cnt_cry_9;
    wire value_cnt_cry_10;
    wire value_cntZ0Z_12;
    wire value_cnt_cry_11_THRU_CO;
    wire value_cnt_cry_11;
    wire value_cntZ0Z_13;
    wire value_cnt_cry_12_THRU_CO;
    wire value_cnt_cry_12;
    wire value_cntZ0Z_14;
    wire value_cnt_cry_13_THRU_CO;
    wire value_cnt_cry_13;
    wire value_cntZ0Z_15;
    wire value_cnt_cry_14_THRU_CO;
    wire value_cnt_cry_14;
    wire value_cnt_cry_15;
    wire value_cntZ0Z_16;
    wire value_cnt_cry_15_THRU_CO;
    wire bfn_6_7_0_;
    wire value_cntZ0Z_17;
    wire value_cnt_cry_16_THRU_CO;
    wire value_cnt_cry_16;
    wire value_cntZ0Z_18;
    wire value_cnt_cry_17_THRU_CO;
    wire value_cnt_cry_17;
    wire value_cntZ0Z_19;
    wire value_cnt_cry_18_THRU_CO;
    wire value_cnt_cry_18;
    wire value_cntZ0Z_20;
    wire value_cnt_cry_19_THRU_CO;
    wire value_cnt_cry_19;
    wire value_cntZ0Z_21;
    wire value_cnt_cry_20_THRU_CO;
    wire value_cnt_cry_20;
    wire value_cntZ0Z_22;
    wire value_cnt_cry_21_THRU_CO;
    wire value_cnt_cry_21;
    wire value_cnt_cry_22;
    wire value_cntZ0Z_23;
    wire leds_c_0;
    wire register10Z0Z_0;
    wire leds_c_1;
    wire leds_c_2;
    wire leds_c_3;
    wire leds_c_4;
    wire leds_c_5;
    wire sl_reg;
    wire register10Z0Z_9;
    wire leds_c_6;
    wire leds_c_7;
    wire un1_sr_reg_0_i;
    wire CONSTANT_ONE_NET;
    wire value_cnt_cry_10_THRU_CO;
    wire value_cntZ0Z_11;
    wire UC_un1_ld_cnt_0_i;
    wire value_cnt_cry_8_THRU_CO;
    wire value_cntZ0Z_9;
    wire _gnd_net_;
    wire clk_c_g;
    wire value_cnte_0_i_g;
    wire reset_c_g;

    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__2702),
            .GLOBALBUFFEROUTPUT(reset_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__2704),
            .DIN(N__2703),
            .DOUT(N__2702),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__2704),
            .PADOUT(N__2703),
            .PADIN(N__2702),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__2692),
            .GLOBALBUFFEROUTPUT(clk_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__2694),
            .DIN(N__2693),
            .DOUT(N__2692),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__2694),
            .PADOUT(N__2693),
            .PADIN(N__2692),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_1_iopad (
            .OE(N__2683),
            .DIN(N__2682),
            .DOUT(N__2681),
            .PACKAGEPIN(leds[1]));
    defparam leds_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_1_preio (
            .PADOEN(N__2683),
            .PADOUT(N__2682),
            .PADIN(N__2681),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1914),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_5_iopad (
            .OE(N__2674),
            .DIN(N__2673),
            .DOUT(N__2672),
            .PACKAGEPIN(leds[5]));
    defparam leds_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_5_preio (
            .PADOEN(N__2674),
            .PADOUT(N__2673),
            .PADIN(N__2672),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2550),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_0_iopad (
            .OE(N__2665),
            .DIN(N__2664),
            .DOUT(N__2663),
            .PACKAGEPIN(leds[0]));
    defparam leds_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_0_preio (
            .PADOEN(N__2665),
            .PADOUT(N__2664),
            .PADIN(N__2663),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1956),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_4_iopad (
            .OE(N__2656),
            .DIN(N__2655),
            .DOUT(N__2654),
            .PACKAGEPIN(leds[4]));
    defparam leds_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_4_preio (
            .PADOEN(N__2656),
            .PADOUT(N__2655),
            .PADIN(N__2654),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2574),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_3_iopad (
            .OE(N__2647),
            .DIN(N__2646),
            .DOUT(N__2645),
            .PACKAGEPIN(leds[3]));
    defparam leds_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_3_preio (
            .PADOEN(N__2647),
            .PADOUT(N__2646),
            .PADIN(N__2645),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2601),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_7_iopad (
            .OE(N__2638),
            .DIN(N__2637),
            .DOUT(N__2636),
            .PACKAGEPIN(leds[7]));
    defparam leds_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_7_preio (
            .PADOEN(N__2638),
            .PADOUT(N__2637),
            .PADIN(N__2636),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2433),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_2_iopad (
            .OE(N__2629),
            .DIN(N__2628),
            .DOUT(N__2627),
            .PACKAGEPIN(leds[2]));
    defparam leds_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_2_preio (
            .PADOEN(N__2629),
            .PADOUT(N__2628),
            .PADIN(N__2627),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1890),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD leds_obuf_6_iopad (
            .OE(N__2620),
            .DIN(N__2619),
            .DOUT(N__2618),
            .PACKAGEPIN(leds[6]));
    defparam leds_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam leds_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO leds_obuf_6_preio (
            .PADOEN(N__2620),
            .PADOUT(N__2619),
            .PADIN(N__2618),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2454),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IoInMux I__598 (
            .O(N__2601),
            .I(N__2598));
    LocalMux I__597 (
            .O(N__2598),
            .I(N__2595));
    IoSpan4Mux I__596 (
            .O(N__2595),
            .I(N__2591));
    CascadeMux I__595 (
            .O(N__2594),
            .I(N__2588));
    Span4Mux_s3_h I__594 (
            .O(N__2591),
            .I(N__2584));
    InMux I__593 (
            .O(N__2588),
            .I(N__2579));
    InMux I__592 (
            .O(N__2587),
            .I(N__2579));
    Odrv4 I__591 (
            .O(N__2584),
            .I(leds_c_3));
    LocalMux I__590 (
            .O(N__2579),
            .I(leds_c_3));
    IoInMux I__589 (
            .O(N__2574),
            .I(N__2571));
    LocalMux I__588 (
            .O(N__2571),
            .I(N__2567));
    CascadeMux I__587 (
            .O(N__2570),
            .I(N__2564));
    Span12Mux_s6_h I__586 (
            .O(N__2567),
            .I(N__2560));
    InMux I__585 (
            .O(N__2564),
            .I(N__2555));
    InMux I__584 (
            .O(N__2563),
            .I(N__2555));
    Odrv12 I__583 (
            .O(N__2560),
            .I(leds_c_4));
    LocalMux I__582 (
            .O(N__2555),
            .I(leds_c_4));
    IoInMux I__581 (
            .O(N__2550),
            .I(N__2547));
    LocalMux I__580 (
            .O(N__2547),
            .I(N__2544));
    Span4Mux_s3_h I__579 (
            .O(N__2544),
            .I(N__2541));
    Span4Mux_v I__578 (
            .O(N__2541),
            .I(N__2536));
    InMux I__577 (
            .O(N__2540),
            .I(N__2531));
    InMux I__576 (
            .O(N__2539),
            .I(N__2531));
    Odrv4 I__575 (
            .O(N__2536),
            .I(leds_c_5));
    LocalMux I__574 (
            .O(N__2531),
            .I(leds_c_5));
    InMux I__573 (
            .O(N__2526),
            .I(N__2505));
    InMux I__572 (
            .O(N__2525),
            .I(N__2505));
    InMux I__571 (
            .O(N__2524),
            .I(N__2505));
    InMux I__570 (
            .O(N__2523),
            .I(N__2505));
    InMux I__569 (
            .O(N__2522),
            .I(N__2505));
    InMux I__568 (
            .O(N__2521),
            .I(N__2505));
    InMux I__567 (
            .O(N__2520),
            .I(N__2505));
    LocalMux I__566 (
            .O(N__2505),
            .I(N__2498));
    InMux I__565 (
            .O(N__2504),
            .I(N__2491));
    InMux I__564 (
            .O(N__2503),
            .I(N__2491));
    InMux I__563 (
            .O(N__2502),
            .I(N__2491));
    InMux I__562 (
            .O(N__2501),
            .I(N__2487));
    Span4Mux_v I__561 (
            .O(N__2498),
            .I(N__2484));
    LocalMux I__560 (
            .O(N__2491),
            .I(N__2481));
    InMux I__559 (
            .O(N__2490),
            .I(N__2478));
    LocalMux I__558 (
            .O(N__2487),
            .I(sl_reg));
    Odrv4 I__557 (
            .O(N__2484),
            .I(sl_reg));
    Odrv4 I__556 (
            .O(N__2481),
            .I(sl_reg));
    LocalMux I__555 (
            .O(N__2478),
            .I(sl_reg));
    InMux I__554 (
            .O(N__2469),
            .I(N__2462));
    InMux I__553 (
            .O(N__2468),
            .I(N__2462));
    InMux I__552 (
            .O(N__2467),
            .I(N__2459));
    LocalMux I__551 (
            .O(N__2462),
            .I(register10Z0Z_9));
    LocalMux I__550 (
            .O(N__2459),
            .I(register10Z0Z_9));
    IoInMux I__549 (
            .O(N__2454),
            .I(N__2451));
    LocalMux I__548 (
            .O(N__2451),
            .I(N__2448));
    Span12Mux_s6_h I__547 (
            .O(N__2448),
            .I(N__2443));
    InMux I__546 (
            .O(N__2447),
            .I(N__2438));
    InMux I__545 (
            .O(N__2446),
            .I(N__2438));
    Odrv12 I__544 (
            .O(N__2443),
            .I(leds_c_6));
    LocalMux I__543 (
            .O(N__2438),
            .I(leds_c_6));
    IoInMux I__542 (
            .O(N__2433),
            .I(N__2430));
    LocalMux I__541 (
            .O(N__2430),
            .I(N__2427));
    IoSpan4Mux I__540 (
            .O(N__2427),
            .I(N__2424));
    Span4Mux_s3_h I__539 (
            .O(N__2424),
            .I(N__2420));
    CascadeMux I__538 (
            .O(N__2423),
            .I(N__2417));
    Span4Mux_v I__537 (
            .O(N__2420),
            .I(N__2413));
    InMux I__536 (
            .O(N__2417),
            .I(N__2408));
    InMux I__535 (
            .O(N__2416),
            .I(N__2408));
    Odrv4 I__534 (
            .O(N__2413),
            .I(leds_c_7));
    LocalMux I__533 (
            .O(N__2408),
            .I(leds_c_7));
    CEMux I__532 (
            .O(N__2403),
            .I(N__2400));
    LocalMux I__531 (
            .O(N__2400),
            .I(N__2397));
    Span4Mux_v I__530 (
            .O(N__2397),
            .I(N__2393));
    CEMux I__529 (
            .O(N__2396),
            .I(N__2390));
    Span4Mux_h I__528 (
            .O(N__2393),
            .I(N__2387));
    LocalMux I__527 (
            .O(N__2390),
            .I(N__2384));
    Odrv4 I__526 (
            .O(N__2387),
            .I(un1_sr_reg_0_i));
    Odrv12 I__525 (
            .O(N__2384),
            .I(un1_sr_reg_0_i));
    CascadeMux I__524 (
            .O(N__2379),
            .I(N__2373));
    InMux I__523 (
            .O(N__2378),
            .I(N__2363));
    InMux I__522 (
            .O(N__2377),
            .I(N__2363));
    InMux I__521 (
            .O(N__2376),
            .I(N__2363));
    InMux I__520 (
            .O(N__2373),
            .I(N__2354));
    InMux I__519 (
            .O(N__2372),
            .I(N__2354));
    InMux I__518 (
            .O(N__2371),
            .I(N__2354));
    InMux I__517 (
            .O(N__2370),
            .I(N__2354));
    LocalMux I__516 (
            .O(N__2363),
            .I(N__2351));
    LocalMux I__515 (
            .O(N__2354),
            .I(N__2333));
    Span4Mux_v I__514 (
            .O(N__2351),
            .I(N__2330));
    InMux I__513 (
            .O(N__2350),
            .I(N__2321));
    InMux I__512 (
            .O(N__2349),
            .I(N__2321));
    InMux I__511 (
            .O(N__2348),
            .I(N__2321));
    InMux I__510 (
            .O(N__2347),
            .I(N__2321));
    InMux I__509 (
            .O(N__2346),
            .I(N__2312));
    InMux I__508 (
            .O(N__2345),
            .I(N__2312));
    InMux I__507 (
            .O(N__2344),
            .I(N__2312));
    InMux I__506 (
            .O(N__2343),
            .I(N__2312));
    InMux I__505 (
            .O(N__2342),
            .I(N__2305));
    InMux I__504 (
            .O(N__2341),
            .I(N__2305));
    InMux I__503 (
            .O(N__2340),
            .I(N__2305));
    InMux I__502 (
            .O(N__2339),
            .I(N__2296));
    InMux I__501 (
            .O(N__2338),
            .I(N__2296));
    InMux I__500 (
            .O(N__2337),
            .I(N__2296));
    InMux I__499 (
            .O(N__2336),
            .I(N__2296));
    Odrv4 I__498 (
            .O(N__2333),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__497 (
            .O(N__2330),
            .I(CONSTANT_ONE_NET));
    LocalMux I__496 (
            .O(N__2321),
            .I(CONSTANT_ONE_NET));
    LocalMux I__495 (
            .O(N__2312),
            .I(CONSTANT_ONE_NET));
    LocalMux I__494 (
            .O(N__2305),
            .I(CONSTANT_ONE_NET));
    LocalMux I__493 (
            .O(N__2296),
            .I(CONSTANT_ONE_NET));
    InMux I__492 (
            .O(N__2283),
            .I(N__2280));
    LocalMux I__491 (
            .O(N__2280),
            .I(value_cnt_cry_10_THRU_CO));
    InMux I__490 (
            .O(N__2277),
            .I(N__2272));
    CascadeMux I__489 (
            .O(N__2276),
            .I(N__2269));
    InMux I__488 (
            .O(N__2275),
            .I(N__2266));
    LocalMux I__487 (
            .O(N__2272),
            .I(N__2263));
    InMux I__486 (
            .O(N__2269),
            .I(N__2260));
    LocalMux I__485 (
            .O(N__2266),
            .I(value_cntZ0Z_11));
    Odrv12 I__484 (
            .O(N__2263),
            .I(value_cntZ0Z_11));
    LocalMux I__483 (
            .O(N__2260),
            .I(value_cntZ0Z_11));
    InMux I__482 (
            .O(N__2253),
            .I(N__2247));
    InMux I__481 (
            .O(N__2252),
            .I(N__2247));
    LocalMux I__480 (
            .O(N__2247),
            .I(N__2230));
    InMux I__479 (
            .O(N__2246),
            .I(N__2215));
    InMux I__478 (
            .O(N__2245),
            .I(N__2215));
    InMux I__477 (
            .O(N__2244),
            .I(N__2215));
    InMux I__476 (
            .O(N__2243),
            .I(N__2215));
    InMux I__475 (
            .O(N__2242),
            .I(N__2215));
    InMux I__474 (
            .O(N__2241),
            .I(N__2215));
    InMux I__473 (
            .O(N__2240),
            .I(N__2215));
    InMux I__472 (
            .O(N__2239),
            .I(N__2199));
    InMux I__471 (
            .O(N__2238),
            .I(N__2199));
    InMux I__470 (
            .O(N__2237),
            .I(N__2199));
    InMux I__469 (
            .O(N__2236),
            .I(N__2199));
    InMux I__468 (
            .O(N__2235),
            .I(N__2199));
    InMux I__467 (
            .O(N__2234),
            .I(N__2199));
    InMux I__466 (
            .O(N__2233),
            .I(N__2199));
    Span4Mux_h I__465 (
            .O(N__2230),
            .I(N__2189));
    LocalMux I__464 (
            .O(N__2215),
            .I(N__2186));
    InMux I__463 (
            .O(N__2214),
            .I(N__2183));
    LocalMux I__462 (
            .O(N__2199),
            .I(N__2180));
    InMux I__461 (
            .O(N__2198),
            .I(N__2175));
    InMux I__460 (
            .O(N__2197),
            .I(N__2175));
    InMux I__459 (
            .O(N__2196),
            .I(N__2164));
    InMux I__458 (
            .O(N__2195),
            .I(N__2164));
    InMux I__457 (
            .O(N__2194),
            .I(N__2164));
    InMux I__456 (
            .O(N__2193),
            .I(N__2164));
    InMux I__455 (
            .O(N__2192),
            .I(N__2164));
    Odrv4 I__454 (
            .O(N__2189),
            .I(UC_un1_ld_cnt_0_i));
    Odrv4 I__453 (
            .O(N__2186),
            .I(UC_un1_ld_cnt_0_i));
    LocalMux I__452 (
            .O(N__2183),
            .I(UC_un1_ld_cnt_0_i));
    Odrv4 I__451 (
            .O(N__2180),
            .I(UC_un1_ld_cnt_0_i));
    LocalMux I__450 (
            .O(N__2175),
            .I(UC_un1_ld_cnt_0_i));
    LocalMux I__449 (
            .O(N__2164),
            .I(UC_un1_ld_cnt_0_i));
    CascadeMux I__448 (
            .O(N__2151),
            .I(N__2148));
    InMux I__447 (
            .O(N__2148),
            .I(N__2145));
    LocalMux I__446 (
            .O(N__2145),
            .I(value_cnt_cry_8_THRU_CO));
    InMux I__445 (
            .O(N__2142),
            .I(N__2137));
    CascadeMux I__444 (
            .O(N__2141),
            .I(N__2134));
    InMux I__443 (
            .O(N__2140),
            .I(N__2131));
    LocalMux I__442 (
            .O(N__2137),
            .I(N__2128));
    InMux I__441 (
            .O(N__2134),
            .I(N__2125));
    LocalMux I__440 (
            .O(N__2131),
            .I(value_cntZ0Z_9));
    Odrv12 I__439 (
            .O(N__2128),
            .I(value_cntZ0Z_9));
    LocalMux I__438 (
            .O(N__2125),
            .I(value_cntZ0Z_9));
    ClkMux I__437 (
            .O(N__2118),
            .I(N__2091));
    ClkMux I__436 (
            .O(N__2117),
            .I(N__2091));
    ClkMux I__435 (
            .O(N__2116),
            .I(N__2091));
    ClkMux I__434 (
            .O(N__2115),
            .I(N__2091));
    ClkMux I__433 (
            .O(N__2114),
            .I(N__2091));
    ClkMux I__432 (
            .O(N__2113),
            .I(N__2091));
    ClkMux I__431 (
            .O(N__2112),
            .I(N__2091));
    ClkMux I__430 (
            .O(N__2111),
            .I(N__2091));
    ClkMux I__429 (
            .O(N__2110),
            .I(N__2091));
    GlobalMux I__428 (
            .O(N__2091),
            .I(N__2088));
    gio2CtrlBuf I__427 (
            .O(N__2088),
            .I(clk_c_g));
    CEMux I__426 (
            .O(N__2085),
            .I(N__2070));
    CEMux I__425 (
            .O(N__2084),
            .I(N__2070));
    CEMux I__424 (
            .O(N__2083),
            .I(N__2070));
    CEMux I__423 (
            .O(N__2082),
            .I(N__2070));
    CEMux I__422 (
            .O(N__2081),
            .I(N__2070));
    GlobalMux I__421 (
            .O(N__2070),
            .I(N__2067));
    gio2CtrlBuf I__420 (
            .O(N__2067),
            .I(value_cnte_0_i_g));
    SRMux I__419 (
            .O(N__2064),
            .I(N__2037));
    SRMux I__418 (
            .O(N__2063),
            .I(N__2037));
    SRMux I__417 (
            .O(N__2062),
            .I(N__2037));
    SRMux I__416 (
            .O(N__2061),
            .I(N__2037));
    SRMux I__415 (
            .O(N__2060),
            .I(N__2037));
    SRMux I__414 (
            .O(N__2059),
            .I(N__2037));
    SRMux I__413 (
            .O(N__2058),
            .I(N__2037));
    SRMux I__412 (
            .O(N__2057),
            .I(N__2037));
    SRMux I__411 (
            .O(N__2056),
            .I(N__2037));
    GlobalMux I__410 (
            .O(N__2037),
            .I(N__2034));
    gio2CtrlBuf I__409 (
            .O(N__2034),
            .I(reset_c_g));
    CascadeMux I__408 (
            .O(N__2031),
            .I(N__2027));
    InMux I__407 (
            .O(N__2030),
            .I(N__2023));
    InMux I__406 (
            .O(N__2027),
            .I(N__2020));
    InMux I__405 (
            .O(N__2026),
            .I(N__2017));
    LocalMux I__404 (
            .O(N__2023),
            .I(value_cntZ0Z_21));
    LocalMux I__403 (
            .O(N__2020),
            .I(value_cntZ0Z_21));
    LocalMux I__402 (
            .O(N__2017),
            .I(value_cntZ0Z_21));
    InMux I__401 (
            .O(N__2010),
            .I(N__2007));
    LocalMux I__400 (
            .O(N__2007),
            .I(value_cnt_cry_20_THRU_CO));
    InMux I__399 (
            .O(N__2004),
            .I(value_cnt_cry_20));
    InMux I__398 (
            .O(N__2001),
            .I(N__1996));
    InMux I__397 (
            .O(N__2000),
            .I(N__1993));
    InMux I__396 (
            .O(N__1999),
            .I(N__1990));
    LocalMux I__395 (
            .O(N__1996),
            .I(value_cntZ0Z_22));
    LocalMux I__394 (
            .O(N__1993),
            .I(value_cntZ0Z_22));
    LocalMux I__393 (
            .O(N__1990),
            .I(value_cntZ0Z_22));
    InMux I__392 (
            .O(N__1983),
            .I(N__1980));
    LocalMux I__391 (
            .O(N__1980),
            .I(value_cnt_cry_21_THRU_CO));
    InMux I__390 (
            .O(N__1977),
            .I(value_cnt_cry_21));
    InMux I__389 (
            .O(N__1974),
            .I(value_cnt_cry_22));
    InMux I__388 (
            .O(N__1971),
            .I(N__1967));
    InMux I__387 (
            .O(N__1970),
            .I(N__1964));
    LocalMux I__386 (
            .O(N__1967),
            .I(N__1961));
    LocalMux I__385 (
            .O(N__1964),
            .I(value_cntZ0Z_23));
    Odrv4 I__384 (
            .O(N__1961),
            .I(value_cntZ0Z_23));
    IoInMux I__383 (
            .O(N__1956),
            .I(N__1953));
    LocalMux I__382 (
            .O(N__1953),
            .I(N__1950));
    Span4Mux_s2_h I__381 (
            .O(N__1950),
            .I(N__1947));
    Span4Mux_h I__380 (
            .O(N__1947),
            .I(N__1942));
    InMux I__379 (
            .O(N__1946),
            .I(N__1937));
    InMux I__378 (
            .O(N__1945),
            .I(N__1937));
    Odrv4 I__377 (
            .O(N__1942),
            .I(leds_c_0));
    LocalMux I__376 (
            .O(N__1937),
            .I(leds_c_0));
    CascadeMux I__375 (
            .O(N__1932),
            .I(N__1929));
    InMux I__374 (
            .O(N__1929),
            .I(N__1922));
    InMux I__373 (
            .O(N__1928),
            .I(N__1922));
    InMux I__372 (
            .O(N__1927),
            .I(N__1919));
    LocalMux I__371 (
            .O(N__1922),
            .I(register10Z0Z_0));
    LocalMux I__370 (
            .O(N__1919),
            .I(register10Z0Z_0));
    IoInMux I__369 (
            .O(N__1914),
            .I(N__1911));
    LocalMux I__368 (
            .O(N__1911),
            .I(N__1908));
    Span12Mux_s6_h I__367 (
            .O(N__1908),
            .I(N__1903));
    InMux I__366 (
            .O(N__1907),
            .I(N__1900));
    InMux I__365 (
            .O(N__1906),
            .I(N__1897));
    Odrv12 I__364 (
            .O(N__1903),
            .I(leds_c_1));
    LocalMux I__363 (
            .O(N__1900),
            .I(leds_c_1));
    LocalMux I__362 (
            .O(N__1897),
            .I(leds_c_1));
    IoInMux I__361 (
            .O(N__1890),
            .I(N__1887));
    LocalMux I__360 (
            .O(N__1887),
            .I(N__1884));
    Span4Mux_s2_h I__359 (
            .O(N__1884),
            .I(N__1881));
    Span4Mux_h I__358 (
            .O(N__1881),
            .I(N__1876));
    InMux I__357 (
            .O(N__1880),
            .I(N__1873));
    InMux I__356 (
            .O(N__1879),
            .I(N__1870));
    Odrv4 I__355 (
            .O(N__1876),
            .I(leds_c_2));
    LocalMux I__354 (
            .O(N__1873),
            .I(leds_c_2));
    LocalMux I__353 (
            .O(N__1870),
            .I(leds_c_2));
    CascadeMux I__352 (
            .O(N__1863),
            .I(N__1858));
    InMux I__351 (
            .O(N__1862),
            .I(N__1855));
    InMux I__350 (
            .O(N__1861),
            .I(N__1852));
    InMux I__349 (
            .O(N__1858),
            .I(N__1849));
    LocalMux I__348 (
            .O(N__1855),
            .I(value_cntZ0Z_13));
    LocalMux I__347 (
            .O(N__1852),
            .I(value_cntZ0Z_13));
    LocalMux I__346 (
            .O(N__1849),
            .I(value_cntZ0Z_13));
    InMux I__345 (
            .O(N__1842),
            .I(N__1839));
    LocalMux I__344 (
            .O(N__1839),
            .I(value_cnt_cry_12_THRU_CO));
    InMux I__343 (
            .O(N__1836),
            .I(value_cnt_cry_12));
    CascadeMux I__342 (
            .O(N__1833),
            .I(N__1828));
    CascadeMux I__341 (
            .O(N__1832),
            .I(N__1825));
    InMux I__340 (
            .O(N__1831),
            .I(N__1822));
    InMux I__339 (
            .O(N__1828),
            .I(N__1819));
    InMux I__338 (
            .O(N__1825),
            .I(N__1816));
    LocalMux I__337 (
            .O(N__1822),
            .I(value_cntZ0Z_14));
    LocalMux I__336 (
            .O(N__1819),
            .I(value_cntZ0Z_14));
    LocalMux I__335 (
            .O(N__1816),
            .I(value_cntZ0Z_14));
    InMux I__334 (
            .O(N__1809),
            .I(N__1806));
    LocalMux I__333 (
            .O(N__1806),
            .I(value_cnt_cry_13_THRU_CO));
    InMux I__332 (
            .O(N__1803),
            .I(value_cnt_cry_13));
    CascadeMux I__331 (
            .O(N__1800),
            .I(N__1795));
    InMux I__330 (
            .O(N__1799),
            .I(N__1792));
    InMux I__329 (
            .O(N__1798),
            .I(N__1789));
    InMux I__328 (
            .O(N__1795),
            .I(N__1786));
    LocalMux I__327 (
            .O(N__1792),
            .I(value_cntZ0Z_15));
    LocalMux I__326 (
            .O(N__1789),
            .I(value_cntZ0Z_15));
    LocalMux I__325 (
            .O(N__1786),
            .I(value_cntZ0Z_15));
    InMux I__324 (
            .O(N__1779),
            .I(N__1776));
    LocalMux I__323 (
            .O(N__1776),
            .I(value_cnt_cry_14_THRU_CO));
    InMux I__322 (
            .O(N__1773),
            .I(value_cnt_cry_14));
    CascadeMux I__321 (
            .O(N__1770),
            .I(N__1765));
    InMux I__320 (
            .O(N__1769),
            .I(N__1762));
    InMux I__319 (
            .O(N__1768),
            .I(N__1759));
    InMux I__318 (
            .O(N__1765),
            .I(N__1756));
    LocalMux I__317 (
            .O(N__1762),
            .I(value_cntZ0Z_16));
    LocalMux I__316 (
            .O(N__1759),
            .I(value_cntZ0Z_16));
    LocalMux I__315 (
            .O(N__1756),
            .I(value_cntZ0Z_16));
    InMux I__314 (
            .O(N__1749),
            .I(N__1746));
    LocalMux I__313 (
            .O(N__1746),
            .I(value_cnt_cry_15_THRU_CO));
    InMux I__312 (
            .O(N__1743),
            .I(bfn_6_7_0_));
    CascadeMux I__311 (
            .O(N__1740),
            .I(N__1736));
    InMux I__310 (
            .O(N__1739),
            .I(N__1732));
    InMux I__309 (
            .O(N__1736),
            .I(N__1729));
    InMux I__308 (
            .O(N__1735),
            .I(N__1726));
    LocalMux I__307 (
            .O(N__1732),
            .I(value_cntZ0Z_17));
    LocalMux I__306 (
            .O(N__1729),
            .I(value_cntZ0Z_17));
    LocalMux I__305 (
            .O(N__1726),
            .I(value_cntZ0Z_17));
    InMux I__304 (
            .O(N__1719),
            .I(N__1716));
    LocalMux I__303 (
            .O(N__1716),
            .I(value_cnt_cry_16_THRU_CO));
    InMux I__302 (
            .O(N__1713),
            .I(value_cnt_cry_16));
    CascadeMux I__301 (
            .O(N__1710),
            .I(N__1705));
    CascadeMux I__300 (
            .O(N__1709),
            .I(N__1702));
    InMux I__299 (
            .O(N__1708),
            .I(N__1699));
    InMux I__298 (
            .O(N__1705),
            .I(N__1696));
    InMux I__297 (
            .O(N__1702),
            .I(N__1693));
    LocalMux I__296 (
            .O(N__1699),
            .I(value_cntZ0Z_18));
    LocalMux I__295 (
            .O(N__1696),
            .I(value_cntZ0Z_18));
    LocalMux I__294 (
            .O(N__1693),
            .I(value_cntZ0Z_18));
    InMux I__293 (
            .O(N__1686),
            .I(N__1683));
    LocalMux I__292 (
            .O(N__1683),
            .I(value_cnt_cry_17_THRU_CO));
    InMux I__291 (
            .O(N__1680),
            .I(value_cnt_cry_17));
    CascadeMux I__290 (
            .O(N__1677),
            .I(N__1673));
    InMux I__289 (
            .O(N__1676),
            .I(N__1669));
    InMux I__288 (
            .O(N__1673),
            .I(N__1666));
    InMux I__287 (
            .O(N__1672),
            .I(N__1663));
    LocalMux I__286 (
            .O(N__1669),
            .I(value_cntZ0Z_19));
    LocalMux I__285 (
            .O(N__1666),
            .I(value_cntZ0Z_19));
    LocalMux I__284 (
            .O(N__1663),
            .I(value_cntZ0Z_19));
    InMux I__283 (
            .O(N__1656),
            .I(N__1653));
    LocalMux I__282 (
            .O(N__1653),
            .I(value_cnt_cry_18_THRU_CO));
    InMux I__281 (
            .O(N__1650),
            .I(value_cnt_cry_18));
    CascadeMux I__280 (
            .O(N__1647),
            .I(N__1642));
    InMux I__279 (
            .O(N__1646),
            .I(N__1639));
    InMux I__278 (
            .O(N__1645),
            .I(N__1636));
    InMux I__277 (
            .O(N__1642),
            .I(N__1633));
    LocalMux I__276 (
            .O(N__1639),
            .I(value_cntZ0Z_20));
    LocalMux I__275 (
            .O(N__1636),
            .I(value_cntZ0Z_20));
    LocalMux I__274 (
            .O(N__1633),
            .I(value_cntZ0Z_20));
    InMux I__273 (
            .O(N__1626),
            .I(N__1623));
    LocalMux I__272 (
            .O(N__1623),
            .I(value_cnt_cry_19_THRU_CO));
    InMux I__271 (
            .O(N__1620),
            .I(value_cnt_cry_19));
    CascadeMux I__270 (
            .O(N__1617),
            .I(N__1612));
    InMux I__269 (
            .O(N__1616),
            .I(N__1609));
    InMux I__268 (
            .O(N__1615),
            .I(N__1606));
    InMux I__267 (
            .O(N__1612),
            .I(N__1603));
    LocalMux I__266 (
            .O(N__1609),
            .I(value_cntZ0Z_5));
    LocalMux I__265 (
            .O(N__1606),
            .I(value_cntZ0Z_5));
    LocalMux I__264 (
            .O(N__1603),
            .I(value_cntZ0Z_5));
    InMux I__263 (
            .O(N__1596),
            .I(N__1593));
    LocalMux I__262 (
            .O(N__1593),
            .I(value_cnt_cry_4_THRU_CO));
    InMux I__261 (
            .O(N__1590),
            .I(value_cnt_cry_4));
    CascadeMux I__260 (
            .O(N__1587),
            .I(N__1582));
    CascadeMux I__259 (
            .O(N__1586),
            .I(N__1579));
    InMux I__258 (
            .O(N__1585),
            .I(N__1576));
    InMux I__257 (
            .O(N__1582),
            .I(N__1573));
    InMux I__256 (
            .O(N__1579),
            .I(N__1570));
    LocalMux I__255 (
            .O(N__1576),
            .I(value_cntZ0Z_6));
    LocalMux I__254 (
            .O(N__1573),
            .I(value_cntZ0Z_6));
    LocalMux I__253 (
            .O(N__1570),
            .I(value_cntZ0Z_6));
    InMux I__252 (
            .O(N__1563),
            .I(N__1560));
    LocalMux I__251 (
            .O(N__1560),
            .I(value_cnt_cry_5_THRU_CO));
    InMux I__250 (
            .O(N__1557),
            .I(value_cnt_cry_5));
    CascadeMux I__249 (
            .O(N__1554),
            .I(N__1549));
    InMux I__248 (
            .O(N__1553),
            .I(N__1546));
    InMux I__247 (
            .O(N__1552),
            .I(N__1543));
    InMux I__246 (
            .O(N__1549),
            .I(N__1540));
    LocalMux I__245 (
            .O(N__1546),
            .I(value_cntZ0Z_7));
    LocalMux I__244 (
            .O(N__1543),
            .I(value_cntZ0Z_7));
    LocalMux I__243 (
            .O(N__1540),
            .I(value_cntZ0Z_7));
    InMux I__242 (
            .O(N__1533),
            .I(N__1530));
    LocalMux I__241 (
            .O(N__1530),
            .I(value_cnt_cry_6_THRU_CO));
    InMux I__240 (
            .O(N__1527),
            .I(value_cnt_cry_6));
    CascadeMux I__239 (
            .O(N__1524),
            .I(N__1519));
    InMux I__238 (
            .O(N__1523),
            .I(N__1516));
    InMux I__237 (
            .O(N__1522),
            .I(N__1513));
    InMux I__236 (
            .O(N__1519),
            .I(N__1510));
    LocalMux I__235 (
            .O(N__1516),
            .I(value_cntZ0Z_8));
    LocalMux I__234 (
            .O(N__1513),
            .I(value_cntZ0Z_8));
    LocalMux I__233 (
            .O(N__1510),
            .I(value_cntZ0Z_8));
    InMux I__232 (
            .O(N__1503),
            .I(N__1500));
    LocalMux I__231 (
            .O(N__1500),
            .I(value_cnt_cry_7_THRU_CO));
    InMux I__230 (
            .O(N__1497),
            .I(bfn_6_6_0_));
    InMux I__229 (
            .O(N__1494),
            .I(value_cnt_cry_8));
    CascadeMux I__228 (
            .O(N__1491),
            .I(N__1486));
    CascadeMux I__227 (
            .O(N__1490),
            .I(N__1483));
    InMux I__226 (
            .O(N__1489),
            .I(N__1480));
    InMux I__225 (
            .O(N__1486),
            .I(N__1477));
    InMux I__224 (
            .O(N__1483),
            .I(N__1474));
    LocalMux I__223 (
            .O(N__1480),
            .I(value_cntZ0Z_10));
    LocalMux I__222 (
            .O(N__1477),
            .I(value_cntZ0Z_10));
    LocalMux I__221 (
            .O(N__1474),
            .I(value_cntZ0Z_10));
    InMux I__220 (
            .O(N__1467),
            .I(N__1464));
    LocalMux I__219 (
            .O(N__1464),
            .I(value_cnt_cry_9_THRU_CO));
    InMux I__218 (
            .O(N__1461),
            .I(value_cnt_cry_9));
    InMux I__217 (
            .O(N__1458),
            .I(value_cnt_cry_10));
    CascadeMux I__216 (
            .O(N__1455),
            .I(N__1450));
    InMux I__215 (
            .O(N__1454),
            .I(N__1447));
    InMux I__214 (
            .O(N__1453),
            .I(N__1444));
    InMux I__213 (
            .O(N__1450),
            .I(N__1441));
    LocalMux I__212 (
            .O(N__1447),
            .I(value_cntZ0Z_12));
    LocalMux I__211 (
            .O(N__1444),
            .I(value_cntZ0Z_12));
    LocalMux I__210 (
            .O(N__1441),
            .I(value_cntZ0Z_12));
    InMux I__209 (
            .O(N__1434),
            .I(N__1431));
    LocalMux I__208 (
            .O(N__1431),
            .I(value_cnt_cry_11_THRU_CO));
    InMux I__207 (
            .O(N__1428),
            .I(value_cnt_cry_11));
    InMux I__206 (
            .O(N__1425),
            .I(N__1419));
    InMux I__205 (
            .O(N__1424),
            .I(N__1419));
    LocalMux I__204 (
            .O(N__1419),
            .I(\UC.epZ0Z_0 ));
    InMux I__203 (
            .O(N__1416),
            .I(N__1413));
    LocalMux I__202 (
            .O(N__1413),
            .I(\UC.epZ0Z_8 ));
    InMux I__201 (
            .O(N__1410),
            .I(N__1404));
    InMux I__200 (
            .O(N__1409),
            .I(N__1404));
    LocalMux I__199 (
            .O(N__1404),
            .I(\UC.epZ0Z_1 ));
    InMux I__198 (
            .O(N__1401),
            .I(N__1396));
    InMux I__197 (
            .O(N__1400),
            .I(N__1393));
    InMux I__196 (
            .O(N__1399),
            .I(N__1390));
    LocalMux I__195 (
            .O(N__1396),
            .I(\UC.epZ0Z_7 ));
    LocalMux I__194 (
            .O(N__1393),
            .I(\UC.epZ0Z_7 ));
    LocalMux I__193 (
            .O(N__1390),
            .I(\UC.epZ0Z_7 ));
    InMux I__192 (
            .O(N__1383),
            .I(N__1378));
    InMux I__191 (
            .O(N__1382),
            .I(N__1375));
    InMux I__190 (
            .O(N__1381),
            .I(N__1372));
    LocalMux I__189 (
            .O(N__1378),
            .I(value_cntZ0Z_0));
    LocalMux I__188 (
            .O(N__1375),
            .I(value_cntZ0Z_0));
    LocalMux I__187 (
            .O(N__1372),
            .I(value_cntZ0Z_0));
    CascadeMux I__186 (
            .O(N__1365),
            .I(N__1360));
    InMux I__185 (
            .O(N__1364),
            .I(N__1357));
    InMux I__184 (
            .O(N__1363),
            .I(N__1354));
    InMux I__183 (
            .O(N__1360),
            .I(N__1351));
    LocalMux I__182 (
            .O(N__1357),
            .I(value_cntZ0Z_1));
    LocalMux I__181 (
            .O(N__1354),
            .I(value_cntZ0Z_1));
    LocalMux I__180 (
            .O(N__1351),
            .I(value_cntZ0Z_1));
    InMux I__179 (
            .O(N__1344),
            .I(N__1341));
    LocalMux I__178 (
            .O(N__1341),
            .I(value_cnt_cry_0_THRU_CO));
    InMux I__177 (
            .O(N__1338),
            .I(value_cnt_cry_0));
    CascadeMux I__176 (
            .O(N__1335),
            .I(N__1330));
    CascadeMux I__175 (
            .O(N__1334),
            .I(N__1327));
    InMux I__174 (
            .O(N__1333),
            .I(N__1324));
    InMux I__173 (
            .O(N__1330),
            .I(N__1321));
    InMux I__172 (
            .O(N__1327),
            .I(N__1318));
    LocalMux I__171 (
            .O(N__1324),
            .I(value_cntZ0Z_2));
    LocalMux I__170 (
            .O(N__1321),
            .I(value_cntZ0Z_2));
    LocalMux I__169 (
            .O(N__1318),
            .I(value_cntZ0Z_2));
    InMux I__168 (
            .O(N__1311),
            .I(N__1308));
    LocalMux I__167 (
            .O(N__1308),
            .I(value_cnt_cry_1_THRU_CO));
    InMux I__166 (
            .O(N__1305),
            .I(value_cnt_cry_1));
    CascadeMux I__165 (
            .O(N__1302),
            .I(N__1297));
    InMux I__164 (
            .O(N__1301),
            .I(N__1294));
    InMux I__163 (
            .O(N__1300),
            .I(N__1291));
    InMux I__162 (
            .O(N__1297),
            .I(N__1288));
    LocalMux I__161 (
            .O(N__1294),
            .I(value_cntZ0Z_3));
    LocalMux I__160 (
            .O(N__1291),
            .I(value_cntZ0Z_3));
    LocalMux I__159 (
            .O(N__1288),
            .I(value_cntZ0Z_3));
    InMux I__158 (
            .O(N__1281),
            .I(N__1278));
    LocalMux I__157 (
            .O(N__1278),
            .I(value_cnt_cry_2_THRU_CO));
    InMux I__156 (
            .O(N__1275),
            .I(value_cnt_cry_2));
    CascadeMux I__155 (
            .O(N__1272),
            .I(N__1267));
    InMux I__154 (
            .O(N__1271),
            .I(N__1264));
    InMux I__153 (
            .O(N__1270),
            .I(N__1261));
    InMux I__152 (
            .O(N__1267),
            .I(N__1258));
    LocalMux I__151 (
            .O(N__1264),
            .I(value_cntZ0Z_4));
    LocalMux I__150 (
            .O(N__1261),
            .I(value_cntZ0Z_4));
    LocalMux I__149 (
            .O(N__1258),
            .I(value_cntZ0Z_4));
    InMux I__148 (
            .O(N__1251),
            .I(N__1248));
    LocalMux I__147 (
            .O(N__1248),
            .I(value_cnt_cry_3_THRU_CO));
    InMux I__146 (
            .O(N__1245),
            .I(value_cnt_cry_3));
    InMux I__145 (
            .O(N__1242),
            .I(N__1237));
    InMux I__144 (
            .O(N__1241),
            .I(N__1234));
    InMux I__143 (
            .O(N__1240),
            .I(N__1231));
    LocalMux I__142 (
            .O(N__1237),
            .I(\UC.epZ0Z_4 ));
    LocalMux I__141 (
            .O(N__1234),
            .I(\UC.epZ0Z_4 ));
    LocalMux I__140 (
            .O(N__1231),
            .I(\UC.epZ0Z_4 ));
    InMux I__139 (
            .O(N__1224),
            .I(N__1220));
    InMux I__138 (
            .O(N__1223),
            .I(N__1217));
    LocalMux I__137 (
            .O(N__1220),
            .I(\UC.sr_reg ));
    LocalMux I__136 (
            .O(N__1217),
            .I(\UC.sr_reg ));
    CascadeMux I__135 (
            .O(N__1212),
            .I(N__1207));
    CascadeMux I__134 (
            .O(N__1211),
            .I(N__1204));
    InMux I__133 (
            .O(N__1210),
            .I(N__1194));
    InMux I__132 (
            .O(N__1207),
            .I(N__1194));
    InMux I__131 (
            .O(N__1204),
            .I(N__1194));
    InMux I__130 (
            .O(N__1203),
            .I(N__1194));
    LocalMux I__129 (
            .O(N__1194),
            .I(op_eq_un4_fin_cnt_20));
    CascadeMux I__128 (
            .O(N__1191),
            .I(N__1186));
    InMux I__127 (
            .O(N__1190),
            .I(N__1180));
    InMux I__126 (
            .O(N__1189),
            .I(N__1180));
    InMux I__125 (
            .O(N__1186),
            .I(N__1175));
    InMux I__124 (
            .O(N__1185),
            .I(N__1175));
    LocalMux I__123 (
            .O(N__1180),
            .I(op_eq_un4_fin_cnt_21));
    LocalMux I__122 (
            .O(N__1175),
            .I(op_eq_un4_fin_cnt_21));
    InMux I__121 (
            .O(N__1170),
            .I(N__1163));
    InMux I__120 (
            .O(N__1169),
            .I(N__1163));
    InMux I__119 (
            .O(N__1168),
            .I(N__1160));
    LocalMux I__118 (
            .O(N__1163),
            .I(\UC.epZ0Z_3 ));
    LocalMux I__117 (
            .O(N__1160),
            .I(\UC.epZ0Z_3 ));
    CascadeMux I__116 (
            .O(N__1155),
            .I(N__1150));
    InMux I__115 (
            .O(N__1154),
            .I(N__1145));
    InMux I__114 (
            .O(N__1153),
            .I(N__1145));
    InMux I__113 (
            .O(N__1150),
            .I(N__1142));
    LocalMux I__112 (
            .O(N__1145),
            .I(\UC.epZ0Z_6 ));
    LocalMux I__111 (
            .O(N__1142),
            .I(\UC.epZ0Z_6 ));
    IoInMux I__110 (
            .O(N__1137),
            .I(N__1134));
    LocalMux I__109 (
            .O(N__1134),
            .I(N__1131));
    Span4Mux_s0_h I__108 (
            .O(N__1131),
            .I(N__1128));
    Odrv4 I__107 (
            .O(N__1128),
            .I(\UC.value_cnte_0_i ));
    CascadeMux I__106 (
            .O(N__1125),
            .I(op_eq_un4_fin_cnt_20_3_cascade_));
    InMux I__105 (
            .O(N__1122),
            .I(N__1119));
    LocalMux I__104 (
            .O(N__1119),
            .I(op_eq_un4_fin_cnt_20_4));
    InMux I__103 (
            .O(N__1116),
            .I(N__1113));
    LocalMux I__102 (
            .O(N__1113),
            .I(op_eq_un4_fin_cnt_21_9));
    InMux I__101 (
            .O(N__1110),
            .I(N__1107));
    LocalMux I__100 (
            .O(N__1107),
            .I(op_eq_un4_fin_cnt_21_11));
    CascadeMux I__99 (
            .O(N__1104),
            .I(N__1101));
    InMux I__98 (
            .O(N__1101),
            .I(N__1098));
    LocalMux I__97 (
            .O(N__1098),
            .I(op_eq_un4_fin_cnt_21_10));
    InMux I__96 (
            .O(N__1095),
            .I(N__1092));
    LocalMux I__95 (
            .O(N__1092),
            .I(op_eq_un4_fin_cnt_21_8));
    defparam IN_MUX_bfv_6_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_5_0_));
    defparam IN_MUX_bfv_6_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_6_0_ (
            .carryinitin(value_cnt_cry_7),
            .carryinitout(bfn_6_6_0_));
    defparam IN_MUX_bfv_6_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_7_0_ (
            .carryinitin(value_cnt_cry_15),
            .carryinitout(bfn_6_7_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB \UC.ep_RNI0P1C_0_3  (
            .USERSIGNALTOGLOBALBUFFER(N__1137),
            .GLOBALBUFFEROUTPUT(value_cnte_0_i_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam value_cnt_RNIOUPL1_8_LC_4_6_1.C_ON=1'b0;
    defparam value_cnt_RNIOUPL1_8_LC_4_6_1.SEQ_MODE=4'b0000;
    defparam value_cnt_RNIOUPL1_8_LC_4_6_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 value_cnt_RNIOUPL1_8_LC_4_6_1 (
            .in0(N__2142),
            .in1(N__1522),
            .in2(N__1491),
            .in3(N__2277),
            .lcout(op_eq_un4_fin_cnt_21_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_RNIMPFN1_12_LC_4_6_2.C_ON=1'b0;
    defparam value_cnt_RNIMPFN1_12_LC_4_6_2.SEQ_MODE=4'b0000;
    defparam value_cnt_RNIMPFN1_12_LC_4_6_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 value_cnt_RNIMPFN1_12_LC_4_6_2 (
            .in0(N__1861),
            .in1(N__1453),
            .in2(N__1833),
            .in3(N__1798),
            .lcout(op_eq_un4_fin_cnt_21_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_RNIQ34K1_4_LC_4_6_4.C_ON=1'b0;
    defparam value_cnt_RNIQ34K1_4_LC_4_6_4.SEQ_MODE=4'b0000;
    defparam value_cnt_RNIQ34K1_4_LC_4_6_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 value_cnt_RNIQ34K1_4_LC_4_6_4 (
            .in0(N__1615),
            .in1(N__1270),
            .in2(N__1587),
            .in3(N__1552),
            .lcout(op_eq_un4_fin_cnt_21_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_RNIAJ3K1_0_LC_4_6_7.C_ON=1'b0;
    defparam value_cnt_RNIAJ3K1_0_LC_4_6_7.SEQ_MODE=4'b0000;
    defparam value_cnt_RNIAJ3K1_0_LC_4_6_7.LUT_INIT=16'b0000000000000001;
    LogicCell40 value_cnt_RNIAJ3K1_0_LC_4_6_7 (
            .in0(N__1363),
            .in1(N__1382),
            .in2(N__1335),
            .in3(N__1300),
            .lcout(op_eq_un4_fin_cnt_21_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_RNI6AGN1_16_LC_4_7_0.C_ON=1'b0;
    defparam value_cnt_RNI6AGN1_16_LC_4_7_0.SEQ_MODE=4'b0000;
    defparam value_cnt_RNI6AGN1_16_LC_4_7_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 value_cnt_RNI6AGN1_16_LC_4_7_0 (
            .in0(N__1735),
            .in1(N__1768),
            .in2(N__1709),
            .in3(N__1672),
            .lcout(op_eq_un4_fin_cnt_20_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_RNINQPR_20_LC_4_7_3.C_ON=1'b0;
    defparam value_cnt_RNINQPR_20_LC_4_7_3.SEQ_MODE=4'b0000;
    defparam value_cnt_RNINQPR_20_LC_4_7_3.LUT_INIT=16'b0000000000110011;
    LogicCell40 value_cnt_RNINQPR_20_LC_4_7_3 (
            .in0(_gnd_net_),
            .in1(N__1645),
            .in2(_gnd_net_),
            .in3(N__2026),
            .lcout(),
            .ltout(op_eq_un4_fin_cnt_20_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_RNIO34F3_23_LC_4_7_4.C_ON=1'b0;
    defparam value_cnt_RNIO34F3_23_LC_4_7_4.SEQ_MODE=4'b0000;
    defparam value_cnt_RNIO34F3_23_LC_4_7_4.LUT_INIT=16'b0001000000000000;
    LogicCell40 value_cnt_RNIO34F3_23_LC_4_7_4 (
            .in0(N__1971),
            .in1(N__1999),
            .in2(N__1125),
            .in3(N__1122),
            .lcout(op_eq_un4_fin_cnt_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_RNIIFHL6_0_LC_4_7_7.C_ON=1'b0;
    defparam value_cnt_RNIIFHL6_0_LC_4_7_7.SEQ_MODE=4'b0000;
    defparam value_cnt_RNIIFHL6_0_LC_4_7_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 value_cnt_RNIIFHL6_0_LC_4_7_7 (
            .in0(N__1116),
            .in1(N__1110),
            .in2(N__1104),
            .in3(N__1095),
            .lcout(op_eq_un4_fin_cnt_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \UC.ep_3_LC_4_8_0 .C_ON=1'b0;
    defparam \UC.ep_3_LC_4_8_0 .SEQ_MODE=4'b1010;
    defparam \UC.ep_3_LC_4_8_0 .LUT_INIT=16'b1111111101001100;
    LogicCell40 \UC.ep_3_LC_4_8_0  (
            .in0(N__1189),
            .in1(N__1169),
            .in2(N__1212),
            .in3(N__1242),
            .lcout(\UC.epZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2110),
            .ce(),
            .sr(N__2063));
    defparam \UC.ep_6_LC_4_8_1 .C_ON=1'b0;
    defparam \UC.ep_6_LC_4_8_1 .SEQ_MODE=4'b1010;
    defparam \UC.ep_6_LC_4_8_1 .LUT_INIT=16'b1100111011101110;
    LogicCell40 \UC.ep_6_LC_4_8_1  (
            .in0(N__1154),
            .in1(N__1401),
            .in2(N__1191),
            .in3(N__1210),
            .lcout(\UC.epZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2110),
            .ce(),
            .sr(N__2063));
    defparam \UC.ep_2_LC_4_8_3 .C_ON=1'b0;
    defparam \UC.ep_2_LC_4_8_3 .SEQ_MODE=4'b1010;
    defparam \UC.ep_2_LC_4_8_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \UC.ep_2_LC_4_8_3  (
            .in0(N__1170),
            .in1(N__1190),
            .in2(_gnd_net_),
            .in3(N__1203),
            .lcout(\UC.sr_reg ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2110),
            .ce(),
            .sr(N__2063));
    defparam \UC.ep_5_LC_4_8_4 .C_ON=1'b0;
    defparam \UC.ep_5_LC_4_8_4 .SEQ_MODE=4'b1010;
    defparam \UC.ep_5_LC_4_8_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \UC.ep_5_LC_4_8_4  (
            .in0(_gnd_net_),
            .in1(N__1153),
            .in2(N__1211),
            .in3(N__1185),
            .lcout(sl_reg),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2110),
            .ce(),
            .sr(N__2063));
    defparam \UC.ep_RNI0P1C_3_LC_4_9_2 .C_ON=1'b0;
    defparam \UC.ep_RNI0P1C_3_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \UC.ep_RNI0P1C_3_LC_4_9_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \UC.ep_RNI0P1C_3_LC_4_9_2  (
            .in0(N__1168),
            .in1(N__1240),
            .in2(N__1155),
            .in3(N__1399),
            .lcout(\UC.value_cnte_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_1_LC_5_5_1.C_ON=1'b0;
    defparam value_cnt_1_LC_5_5_1.SEQ_MODE=4'b1010;
    defparam value_cnt_1_LC_5_5_1.LUT_INIT=16'b0010001000010001;
    LogicCell40 value_cnt_1_LC_5_5_1 (
            .in0(N__1364),
            .in1(N__2240),
            .in2(_gnd_net_),
            .in3(N__1344),
            .lcout(value_cntZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2117),
            .ce(N__2084),
            .sr(N__2056));
    defparam value_cnt_6_LC_5_5_2.C_ON=1'b0;
    defparam value_cnt_6_LC_5_5_2.SEQ_MODE=4'b1010;
    defparam value_cnt_6_LC_5_5_2.LUT_INIT=16'b0100010000010001;
    LogicCell40 value_cnt_6_LC_5_5_2 (
            .in0(N__2245),
            .in1(N__1585),
            .in2(_gnd_net_),
            .in3(N__1563),
            .lcout(value_cntZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2117),
            .ce(N__2084),
            .sr(N__2056));
    defparam value_cnt_7_LC_5_5_3.C_ON=1'b0;
    defparam value_cnt_7_LC_5_5_3.SEQ_MODE=4'b1010;
    defparam value_cnt_7_LC_5_5_3.LUT_INIT=16'b0010001000010001;
    LogicCell40 value_cnt_7_LC_5_5_3 (
            .in0(N__1553),
            .in1(N__2246),
            .in2(_gnd_net_),
            .in3(N__1533),
            .lcout(value_cntZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2117),
            .ce(N__2084),
            .sr(N__2056));
    defparam value_cnt_4_LC_5_5_4.C_ON=1'b0;
    defparam value_cnt_4_LC_5_5_4.SEQ_MODE=4'b1010;
    defparam value_cnt_4_LC_5_5_4.LUT_INIT=16'b0100010000010001;
    LogicCell40 value_cnt_4_LC_5_5_4 (
            .in0(N__2243),
            .in1(N__1271),
            .in2(_gnd_net_),
            .in3(N__1251),
            .lcout(value_cntZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2117),
            .ce(N__2084),
            .sr(N__2056));
    defparam value_cnt_3_LC_5_5_5.C_ON=1'b0;
    defparam value_cnt_3_LC_5_5_5.SEQ_MODE=4'b1010;
    defparam value_cnt_3_LC_5_5_5.LUT_INIT=16'b0010001000010001;
    LogicCell40 value_cnt_3_LC_5_5_5 (
            .in0(N__1301),
            .in1(N__2242),
            .in2(_gnd_net_),
            .in3(N__1281),
            .lcout(value_cntZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2117),
            .ce(N__2084),
            .sr(N__2056));
    defparam value_cnt_2_LC_5_5_6.C_ON=1'b0;
    defparam value_cnt_2_LC_5_5_6.SEQ_MODE=4'b1010;
    defparam value_cnt_2_LC_5_5_6.LUT_INIT=16'b0100010000010001;
    LogicCell40 value_cnt_2_LC_5_5_6 (
            .in0(N__2241),
            .in1(N__1333),
            .in2(_gnd_net_),
            .in3(N__1311),
            .lcout(value_cntZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2117),
            .ce(N__2084),
            .sr(N__2056));
    defparam value_cnt_5_LC_5_5_7.C_ON=1'b0;
    defparam value_cnt_5_LC_5_5_7.SEQ_MODE=4'b1010;
    defparam value_cnt_5_LC_5_5_7.LUT_INIT=16'b0010001000010001;
    LogicCell40 value_cnt_5_LC_5_5_7 (
            .in0(N__1616),
            .in1(N__2244),
            .in2(_gnd_net_),
            .in3(N__1596),
            .lcout(value_cntZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2117),
            .ce(N__2084),
            .sr(N__2056));
    defparam value_cnt_14_LC_5_6_0.C_ON=1'b0;
    defparam value_cnt_14_LC_5_6_0.SEQ_MODE=4'b1010;
    defparam value_cnt_14_LC_5_6_0.LUT_INIT=16'b0100010000010001;
    LogicCell40 value_cnt_14_LC_5_6_0 (
            .in0(N__2237),
            .in1(N__1831),
            .in2(_gnd_net_),
            .in3(N__1809),
            .lcout(value_cntZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2114),
            .ce(N__2082),
            .sr(N__2058));
    defparam value_cnt_10_LC_5_6_2.C_ON=1'b0;
    defparam value_cnt_10_LC_5_6_2.SEQ_MODE=4'b1010;
    defparam value_cnt_10_LC_5_6_2.LUT_INIT=16'b0100010000010001;
    LogicCell40 value_cnt_10_LC_5_6_2 (
            .in0(N__2234),
            .in1(N__1489),
            .in2(_gnd_net_),
            .in3(N__1467),
            .lcout(value_cntZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2114),
            .ce(N__2082),
            .sr(N__2058));
    defparam value_cnt_0_LC_5_6_3.C_ON=1'b0;
    defparam value_cnt_0_LC_5_6_3.SEQ_MODE=4'b1010;
    defparam value_cnt_0_LC_5_6_3.LUT_INIT=16'b0010001000010001;
    LogicCell40 value_cnt_0_LC_5_6_3 (
            .in0(_gnd_net_),
            .in1(N__2233),
            .in2(_gnd_net_),
            .in3(N__1383),
            .lcout(value_cntZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2114),
            .ce(N__2082),
            .sr(N__2058));
    defparam value_cnt_8_LC_5_6_4.C_ON=1'b0;
    defparam value_cnt_8_LC_5_6_4.SEQ_MODE=4'b1011;
    defparam value_cnt_8_LC_5_6_4.LUT_INIT=16'b1110111010111011;
    LogicCell40 value_cnt_8_LC_5_6_4 (
            .in0(N__2239),
            .in1(N__1523),
            .in2(_gnd_net_),
            .in3(N__1503),
            .lcout(value_cntZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2114),
            .ce(N__2082),
            .sr(N__2058));
    defparam value_cnt_13_LC_5_6_5.C_ON=1'b0;
    defparam value_cnt_13_LC_5_6_5.SEQ_MODE=4'b1010;
    defparam value_cnt_13_LC_5_6_5.LUT_INIT=16'b0010001000010001;
    LogicCell40 value_cnt_13_LC_5_6_5 (
            .in0(N__1862),
            .in1(N__2236),
            .in2(_gnd_net_),
            .in3(N__1842),
            .lcout(value_cntZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2114),
            .ce(N__2082),
            .sr(N__2058));
    defparam value_cnt_12_LC_5_6_6.C_ON=1'b0;
    defparam value_cnt_12_LC_5_6_6.SEQ_MODE=4'b1011;
    defparam value_cnt_12_LC_5_6_6.LUT_INIT=16'b1110111010111011;
    LogicCell40 value_cnt_12_LC_5_6_6 (
            .in0(N__2235),
            .in1(N__1454),
            .in2(_gnd_net_),
            .in3(N__1434),
            .lcout(value_cntZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2114),
            .ce(N__2082),
            .sr(N__2058));
    defparam value_cnt_15_LC_5_6_7.C_ON=1'b0;
    defparam value_cnt_15_LC_5_6_7.SEQ_MODE=4'b1010;
    defparam value_cnt_15_LC_5_6_7.LUT_INIT=16'b0010001000010001;
    LogicCell40 value_cnt_15_LC_5_6_7 (
            .in0(N__1799),
            .in1(N__2238),
            .in2(_gnd_net_),
            .in3(N__1779),
            .lcout(value_cntZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2114),
            .ce(N__2082),
            .sr(N__2058));
    defparam value_cnt_18_LC_5_7_0.C_ON=1'b0;
    defparam value_cnt_18_LC_5_7_0.SEQ_MODE=4'b1011;
    defparam value_cnt_18_LC_5_7_0.LUT_INIT=16'b1110111010111011;
    LogicCell40 value_cnt_18_LC_5_7_0 (
            .in0(N__2193),
            .in1(N__1708),
            .in2(_gnd_net_),
            .in3(N__1686),
            .lcout(value_cntZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2112),
            .ce(N__2081),
            .sr(N__2061));
    defparam value_cnt_22_LC_5_7_1.C_ON=1'b0;
    defparam value_cnt_22_LC_5_7_1.SEQ_MODE=4'b1010;
    defparam value_cnt_22_LC_5_7_1.LUT_INIT=16'b0010001000010001;
    LogicCell40 value_cnt_22_LC_5_7_1 (
            .in0(N__2001),
            .in1(N__2196),
            .in2(_gnd_net_),
            .in3(N__1983),
            .lcout(value_cntZ0Z_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2112),
            .ce(N__2081),
            .sr(N__2061));
    defparam value_cnt_19_LC_5_7_2.C_ON=1'b0;
    defparam value_cnt_19_LC_5_7_2.SEQ_MODE=4'b1010;
    defparam value_cnt_19_LC_5_7_2.LUT_INIT=16'b0100010000010001;
    LogicCell40 value_cnt_19_LC_5_7_2 (
            .in0(N__2194),
            .in1(N__1676),
            .in2(_gnd_net_),
            .in3(N__1656),
            .lcout(value_cntZ0Z_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2112),
            .ce(N__2081),
            .sr(N__2061));
    defparam value_cnt_20_LC_5_7_4.C_ON=1'b0;
    defparam value_cnt_20_LC_5_7_4.SEQ_MODE=4'b1011;
    defparam value_cnt_20_LC_5_7_4.LUT_INIT=16'b1110111010111011;
    LogicCell40 value_cnt_20_LC_5_7_4 (
            .in0(N__2195),
            .in1(N__1646),
            .in2(_gnd_net_),
            .in3(N__1626),
            .lcout(value_cntZ0Z_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2112),
            .ce(N__2081),
            .sr(N__2061));
    defparam value_cnt_17_LC_5_7_5.C_ON=1'b0;
    defparam value_cnt_17_LC_5_7_5.SEQ_MODE=4'b1011;
    defparam value_cnt_17_LC_5_7_5.LUT_INIT=16'b1110111010111011;
    LogicCell40 value_cnt_17_LC_5_7_5 (
            .in0(N__2197),
            .in1(N__1739),
            .in2(_gnd_net_),
            .in3(N__1719),
            .lcout(value_cntZ0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2112),
            .ce(N__2081),
            .sr(N__2061));
    defparam value_cnt_16_LC_5_7_6.C_ON=1'b0;
    defparam value_cnt_16_LC_5_7_6.SEQ_MODE=4'b1011;
    defparam value_cnt_16_LC_5_7_6.LUT_INIT=16'b1110111010111011;
    LogicCell40 value_cnt_16_LC_5_7_6 (
            .in0(N__2192),
            .in1(N__1769),
            .in2(_gnd_net_),
            .in3(N__1749),
            .lcout(value_cntZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2112),
            .ce(N__2081),
            .sr(N__2061));
    defparam value_cnt_21_LC_5_7_7.C_ON=1'b0;
    defparam value_cnt_21_LC_5_7_7.SEQ_MODE=4'b1011;
    defparam value_cnt_21_LC_5_7_7.LUT_INIT=16'b1110111010111011;
    LogicCell40 value_cnt_21_LC_5_7_7 (
            .in0(N__2198),
            .in1(N__2030),
            .in2(_gnd_net_),
            .in3(N__2010),
            .lcout(value_cntZ0Z_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2112),
            .ce(N__2081),
            .sr(N__2061));
    defparam \UC.ep_RNIHT06_4_LC_5_8_1 .C_ON=1'b0;
    defparam \UC.ep_RNIHT06_4_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \UC.ep_RNIHT06_4_LC_5_8_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \UC.ep_RNIHT06_4_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(N__1400),
            .in2(_gnd_net_),
            .in3(N__1241),
            .lcout(UC_un1_ld_cnt_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \UC.ep_RNIDP06_2_LC_5_8_4 .C_ON=1'b0;
    defparam \UC.ep_RNIDP06_2_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \UC.ep_RNIDP06_2_LC_5_8_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \UC.ep_RNIDP06_2_LC_5_8_4  (
            .in0(_gnd_net_),
            .in1(N__1223),
            .in2(_gnd_net_),
            .in3(N__2490),
            .lcout(un1_sr_reg_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \UC.ep_4_LC_5_9_1 .C_ON=1'b0;
    defparam \UC.ep_4_LC_5_9_1 .SEQ_MODE=4'b1010;
    defparam \UC.ep_4_LC_5_9_1 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \UC.ep_4_LC_5_9_1  (
            .in0(N__2469),
            .in1(N__1424),
            .in2(N__1932),
            .in3(N__1410),
            .lcout(\UC.epZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2113),
            .ce(),
            .sr(N__2064));
    defparam \UC.ep_0_LC_5_9_3 .C_ON=1'b0;
    defparam \UC.ep_0_LC_5_9_3 .SEQ_MODE=4'b1010;
    defparam \UC.ep_0_LC_5_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \UC.ep_0_LC_5_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1224),
            .lcout(\UC.epZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2113),
            .ce(),
            .sr(N__2064));
    defparam \UC.ep_8_LC_5_9_4 .C_ON=1'b0;
    defparam \UC.ep_8_LC_5_9_4 .SEQ_MODE=4'b1011;
    defparam \UC.ep_8_LC_5_9_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \UC.ep_8_LC_5_9_4  (
            .in0(N__1425),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1928),
            .lcout(\UC.epZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2113),
            .ce(),
            .sr(N__2064));
    defparam \UC.ep_1_LC_5_9_6 .C_ON=1'b0;
    defparam \UC.ep_1_LC_5_9_6 .SEQ_MODE=4'b1010;
    defparam \UC.ep_1_LC_5_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \UC.ep_1_LC_5_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2501),
            .lcout(\UC.epZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2113),
            .ce(),
            .sr(N__2064));
    defparam \UC.ep_7_LC_5_9_7 .C_ON=1'b0;
    defparam \UC.ep_7_LC_5_9_7 .SEQ_MODE=4'b1010;
    defparam \UC.ep_7_LC_5_9_7 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \UC.ep_7_LC_5_9_7  (
            .in0(N__2468),
            .in1(N__1416),
            .in2(_gnd_net_),
            .in3(N__1409),
            .lcout(\UC.epZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2113),
            .ce(),
            .sr(N__2064));
    defparam value_cnt_cry_c_0_LC_6_5_0.C_ON=1'b1;
    defparam value_cnt_cry_c_0_LC_6_5_0.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_c_0_LC_6_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 value_cnt_cry_c_0_LC_6_5_0 (
            .in0(_gnd_net_),
            .in1(N__1381),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_5_0_),
            .carryout(value_cnt_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_0_THRU_LUT4_0_LC_6_5_1.C_ON=1'b1;
    defparam value_cnt_cry_0_THRU_LUT4_0_LC_6_5_1.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_0_THRU_LUT4_0_LC_6_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_0_THRU_LUT4_0_LC_6_5_1 (
            .in0(_gnd_net_),
            .in1(N__2336),
            .in2(N__1365),
            .in3(N__1338),
            .lcout(value_cnt_cry_0_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_0),
            .carryout(value_cnt_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_1_THRU_LUT4_0_LC_6_5_2.C_ON=1'b1;
    defparam value_cnt_cry_1_THRU_LUT4_0_LC_6_5_2.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_1_THRU_LUT4_0_LC_6_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_1_THRU_LUT4_0_LC_6_5_2 (
            .in0(_gnd_net_),
            .in1(N__2340),
            .in2(N__1334),
            .in3(N__1305),
            .lcout(value_cnt_cry_1_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_1),
            .carryout(value_cnt_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_2_THRU_LUT4_0_LC_6_5_3.C_ON=1'b1;
    defparam value_cnt_cry_2_THRU_LUT4_0_LC_6_5_3.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_2_THRU_LUT4_0_LC_6_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_2_THRU_LUT4_0_LC_6_5_3 (
            .in0(_gnd_net_),
            .in1(N__2337),
            .in2(N__1302),
            .in3(N__1275),
            .lcout(value_cnt_cry_2_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_2),
            .carryout(value_cnt_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_3_THRU_LUT4_0_LC_6_5_4.C_ON=1'b1;
    defparam value_cnt_cry_3_THRU_LUT4_0_LC_6_5_4.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_3_THRU_LUT4_0_LC_6_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_3_THRU_LUT4_0_LC_6_5_4 (
            .in0(_gnd_net_),
            .in1(N__2341),
            .in2(N__1272),
            .in3(N__1245),
            .lcout(value_cnt_cry_3_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_3),
            .carryout(value_cnt_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_4_THRU_LUT4_0_LC_6_5_5.C_ON=1'b1;
    defparam value_cnt_cry_4_THRU_LUT4_0_LC_6_5_5.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_4_THRU_LUT4_0_LC_6_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_4_THRU_LUT4_0_LC_6_5_5 (
            .in0(_gnd_net_),
            .in1(N__2338),
            .in2(N__1617),
            .in3(N__1590),
            .lcout(value_cnt_cry_4_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_4),
            .carryout(value_cnt_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_5_THRU_LUT4_0_LC_6_5_6.C_ON=1'b1;
    defparam value_cnt_cry_5_THRU_LUT4_0_LC_6_5_6.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_5_THRU_LUT4_0_LC_6_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_5_THRU_LUT4_0_LC_6_5_6 (
            .in0(_gnd_net_),
            .in1(N__2342),
            .in2(N__1586),
            .in3(N__1557),
            .lcout(value_cnt_cry_5_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_5),
            .carryout(value_cnt_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_6_THRU_LUT4_0_LC_6_5_7.C_ON=1'b1;
    defparam value_cnt_cry_6_THRU_LUT4_0_LC_6_5_7.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_6_THRU_LUT4_0_LC_6_5_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_6_THRU_LUT4_0_LC_6_5_7 (
            .in0(_gnd_net_),
            .in1(N__2339),
            .in2(N__1554),
            .in3(N__1527),
            .lcout(value_cnt_cry_6_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_6),
            .carryout(value_cnt_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_7_THRU_LUT4_0_LC_6_6_0.C_ON=1'b1;
    defparam value_cnt_cry_7_THRU_LUT4_0_LC_6_6_0.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_7_THRU_LUT4_0_LC_6_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_7_THRU_LUT4_0_LC_6_6_0 (
            .in0(_gnd_net_),
            .in1(N__2349),
            .in2(N__1524),
            .in3(N__1497),
            .lcout(value_cnt_cry_7_THRU_CO),
            .ltout(),
            .carryin(bfn_6_6_0_),
            .carryout(value_cnt_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_8_THRU_LUT4_0_LC_6_6_1.C_ON=1'b1;
    defparam value_cnt_cry_8_THRU_LUT4_0_LC_6_6_1.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_8_THRU_LUT4_0_LC_6_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_8_THRU_LUT4_0_LC_6_6_1 (
            .in0(_gnd_net_),
            .in1(N__2346),
            .in2(N__2141),
            .in3(N__1494),
            .lcout(value_cnt_cry_8_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_8),
            .carryout(value_cnt_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_9_THRU_LUT4_0_LC_6_6_2.C_ON=1'b1;
    defparam value_cnt_cry_9_THRU_LUT4_0_LC_6_6_2.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_9_THRU_LUT4_0_LC_6_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_9_THRU_LUT4_0_LC_6_6_2 (
            .in0(_gnd_net_),
            .in1(N__2350),
            .in2(N__1490),
            .in3(N__1461),
            .lcout(value_cnt_cry_9_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_9),
            .carryout(value_cnt_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_10_THRU_LUT4_0_LC_6_6_3.C_ON=1'b1;
    defparam value_cnt_cry_10_THRU_LUT4_0_LC_6_6_3.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_10_THRU_LUT4_0_LC_6_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_10_THRU_LUT4_0_LC_6_6_3 (
            .in0(_gnd_net_),
            .in1(N__2343),
            .in2(N__2276),
            .in3(N__1458),
            .lcout(value_cnt_cry_10_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_10),
            .carryout(value_cnt_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_11_THRU_LUT4_0_LC_6_6_4.C_ON=1'b1;
    defparam value_cnt_cry_11_THRU_LUT4_0_LC_6_6_4.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_11_THRU_LUT4_0_LC_6_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_11_THRU_LUT4_0_LC_6_6_4 (
            .in0(_gnd_net_),
            .in1(N__2347),
            .in2(N__1455),
            .in3(N__1428),
            .lcout(value_cnt_cry_11_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_11),
            .carryout(value_cnt_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_12_THRU_LUT4_0_LC_6_6_5.C_ON=1'b1;
    defparam value_cnt_cry_12_THRU_LUT4_0_LC_6_6_5.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_12_THRU_LUT4_0_LC_6_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_12_THRU_LUT4_0_LC_6_6_5 (
            .in0(_gnd_net_),
            .in1(N__2344),
            .in2(N__1863),
            .in3(N__1836),
            .lcout(value_cnt_cry_12_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_12),
            .carryout(value_cnt_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_13_THRU_LUT4_0_LC_6_6_6.C_ON=1'b1;
    defparam value_cnt_cry_13_THRU_LUT4_0_LC_6_6_6.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_13_THRU_LUT4_0_LC_6_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_13_THRU_LUT4_0_LC_6_6_6 (
            .in0(_gnd_net_),
            .in1(N__2348),
            .in2(N__1832),
            .in3(N__1803),
            .lcout(value_cnt_cry_13_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_13),
            .carryout(value_cnt_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_14_THRU_LUT4_0_LC_6_6_7.C_ON=1'b1;
    defparam value_cnt_cry_14_THRU_LUT4_0_LC_6_6_7.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_14_THRU_LUT4_0_LC_6_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_14_THRU_LUT4_0_LC_6_6_7 (
            .in0(_gnd_net_),
            .in1(N__2345),
            .in2(N__1800),
            .in3(N__1773),
            .lcout(value_cnt_cry_14_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_14),
            .carryout(value_cnt_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_15_THRU_LUT4_0_LC_6_7_0.C_ON=1'b1;
    defparam value_cnt_cry_15_THRU_LUT4_0_LC_6_7_0.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_15_THRU_LUT4_0_LC_6_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_15_THRU_LUT4_0_LC_6_7_0 (
            .in0(_gnd_net_),
            .in1(N__2376),
            .in2(N__1770),
            .in3(N__1743),
            .lcout(value_cnt_cry_15_THRU_CO),
            .ltout(),
            .carryin(bfn_6_7_0_),
            .carryout(value_cnt_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_16_THRU_LUT4_0_LC_6_7_1.C_ON=1'b1;
    defparam value_cnt_cry_16_THRU_LUT4_0_LC_6_7_1.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_16_THRU_LUT4_0_LC_6_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_16_THRU_LUT4_0_LC_6_7_1 (
            .in0(_gnd_net_),
            .in1(N__2370),
            .in2(N__1740),
            .in3(N__1713),
            .lcout(value_cnt_cry_16_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_16),
            .carryout(value_cnt_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_17_THRU_LUT4_0_LC_6_7_2.C_ON=1'b1;
    defparam value_cnt_cry_17_THRU_LUT4_0_LC_6_7_2.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_17_THRU_LUT4_0_LC_6_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_17_THRU_LUT4_0_LC_6_7_2 (
            .in0(_gnd_net_),
            .in1(N__2377),
            .in2(N__1710),
            .in3(N__1680),
            .lcout(value_cnt_cry_17_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_17),
            .carryout(value_cnt_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_18_THRU_LUT4_0_LC_6_7_3.C_ON=1'b1;
    defparam value_cnt_cry_18_THRU_LUT4_0_LC_6_7_3.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_18_THRU_LUT4_0_LC_6_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_18_THRU_LUT4_0_LC_6_7_3 (
            .in0(_gnd_net_),
            .in1(N__2371),
            .in2(N__1677),
            .in3(N__1650),
            .lcout(value_cnt_cry_18_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_18),
            .carryout(value_cnt_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_19_THRU_LUT4_0_LC_6_7_4.C_ON=1'b1;
    defparam value_cnt_cry_19_THRU_LUT4_0_LC_6_7_4.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_19_THRU_LUT4_0_LC_6_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_19_THRU_LUT4_0_LC_6_7_4 (
            .in0(_gnd_net_),
            .in1(N__2378),
            .in2(N__1647),
            .in3(N__1620),
            .lcout(value_cnt_cry_19_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_19),
            .carryout(value_cnt_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_20_THRU_LUT4_0_LC_6_7_5.C_ON=1'b1;
    defparam value_cnt_cry_20_THRU_LUT4_0_LC_6_7_5.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_20_THRU_LUT4_0_LC_6_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_20_THRU_LUT4_0_LC_6_7_5 (
            .in0(_gnd_net_),
            .in1(N__2372),
            .in2(N__2031),
            .in3(N__2004),
            .lcout(value_cnt_cry_20_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_20),
            .carryout(value_cnt_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_cry_21_THRU_LUT4_0_LC_6_7_6.C_ON=1'b1;
    defparam value_cnt_cry_21_THRU_LUT4_0_LC_6_7_6.SEQ_MODE=4'b0000;
    defparam value_cnt_cry_21_THRU_LUT4_0_LC_6_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 value_cnt_cry_21_THRU_LUT4_0_LC_6_7_6 (
            .in0(_gnd_net_),
            .in1(N__2000),
            .in2(N__2379),
            .in3(N__1977),
            .lcout(value_cnt_cry_21_THRU_CO),
            .ltout(),
            .carryin(value_cnt_cry_21),
            .carryout(value_cnt_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_23_LC_6_7_7.C_ON=1'b0;
    defparam value_cnt_23_LC_6_7_7.SEQ_MODE=4'b1011;
    defparam value_cnt_23_LC_6_7_7.LUT_INIT=16'b1110111011011101;
    LogicCell40 value_cnt_23_LC_6_7_7 (
            .in0(N__1970),
            .in1(N__2214),
            .in2(_gnd_net_),
            .in3(N__1974),
            .lcout(value_cntZ0Z_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2115),
            .ce(N__2083),
            .sr(N__2057));
    defparam register10_1_LC_6_8_0.C_ON=1'b0;
    defparam register10_1_LC_6_8_0.SEQ_MODE=4'b1010;
    defparam register10_1_LC_6_8_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 register10_1_LC_6_8_0 (
            .in0(N__2503),
            .in1(N__1927),
            .in2(_gnd_net_),
            .in3(N__1906),
            .lcout(leds_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2111),
            .ce(N__2396),
            .sr(N__2060));
    defparam register10_2_LC_6_8_3.C_ON=1'b0;
    defparam register10_2_LC_6_8_3.SEQ_MODE=4'b1010;
    defparam register10_2_LC_6_8_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 register10_2_LC_6_8_3 (
            .in0(N__1946),
            .in1(N__1880),
            .in2(_gnd_net_),
            .in3(N__2504),
            .lcout(leds_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2111),
            .ce(N__2396),
            .sr(N__2060));
    defparam register10_0_LC_6_8_5.C_ON=1'b0;
    defparam register10_0_LC_6_8_5.SEQ_MODE=4'b1011;
    defparam register10_0_LC_6_8_5.LUT_INIT=16'b0000000010101010;
    LogicCell40 register10_0_LC_6_8_5 (
            .in0(N__1945),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2502),
            .lcout(register10Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2111),
            .ce(N__2396),
            .sr(N__2060));
    defparam register10_3_LC_6_9_0.C_ON=1'b0;
    defparam register10_3_LC_6_9_0.SEQ_MODE=4'b1010;
    defparam register10_3_LC_6_9_0.LUT_INIT=16'b1111101001010000;
    LogicCell40 register10_3_LC_6_9_0 (
            .in0(N__2521),
            .in1(_gnd_net_),
            .in2(N__2594),
            .in3(N__1907),
            .lcout(leds_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2116),
            .ce(N__2403),
            .sr(N__2062));
    defparam register10_6_LC_6_9_1.C_ON=1'b0;
    defparam register10_6_LC_6_9_1.SEQ_MODE=4'b1010;
    defparam register10_6_LC_6_9_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 register10_6_LC_6_9_1 (
            .in0(N__2447),
            .in1(N__2563),
            .in2(_gnd_net_),
            .in3(N__2524),
            .lcout(leds_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2116),
            .ce(N__2403),
            .sr(N__2062));
    defparam register10_4_LC_6_9_2.C_ON=1'b0;
    defparam register10_4_LC_6_9_2.SEQ_MODE=4'b1010;
    defparam register10_4_LC_6_9_2.LUT_INIT=16'b1111101001010000;
    LogicCell40 register10_4_LC_6_9_2 (
            .in0(N__2522),
            .in1(_gnd_net_),
            .in2(N__2570),
            .in3(N__1879),
            .lcout(leds_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2116),
            .ce(N__2403),
            .sr(N__2062));
    defparam register10_5_LC_6_9_3.C_ON=1'b0;
    defparam register10_5_LC_6_9_3.SEQ_MODE=4'b1010;
    defparam register10_5_LC_6_9_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 register10_5_LC_6_9_3 (
            .in0(N__2540),
            .in1(N__2587),
            .in2(_gnd_net_),
            .in3(N__2523),
            .lcout(leds_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2116),
            .ce(N__2403),
            .sr(N__2062));
    defparam register10_7_LC_6_9_4.C_ON=1'b0;
    defparam register10_7_LC_6_9_4.SEQ_MODE=4'b1010;
    defparam register10_7_LC_6_9_4.LUT_INIT=16'b1111101001010000;
    LogicCell40 register10_7_LC_6_9_4 (
            .in0(N__2525),
            .in1(_gnd_net_),
            .in2(N__2423),
            .in3(N__2539),
            .lcout(leds_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2116),
            .ce(N__2403),
            .sr(N__2062));
    defparam register10_9_LC_6_9_5.C_ON=1'b0;
    defparam register10_9_LC_6_9_5.SEQ_MODE=4'b1010;
    defparam register10_9_LC_6_9_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 register10_9_LC_6_9_5 (
            .in0(_gnd_net_),
            .in1(N__2416),
            .in2(_gnd_net_),
            .in3(N__2520),
            .lcout(register10Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2116),
            .ce(N__2403),
            .sr(N__2062));
    defparam register10_8_LC_6_9_6.C_ON=1'b0;
    defparam register10_8_LC_6_9_6.SEQ_MODE=4'b1010;
    defparam register10_8_LC_6_9_6.LUT_INIT=16'b1110111001000100;
    LogicCell40 register10_8_LC_6_9_6 (
            .in0(N__2526),
            .in1(N__2467),
            .in2(_gnd_net_),
            .in3(N__2446),
            .lcout(leds_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2116),
            .ce(N__2403),
            .sr(N__2062));
    defparam CONSTANT_ONE_LUT4_LC_7_5_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_7_5_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_7_5_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_7_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam value_cnt_11_LC_7_6_0.C_ON=1'b0;
    defparam value_cnt_11_LC_7_6_0.SEQ_MODE=4'b1011;
    defparam value_cnt_11_LC_7_6_0.LUT_INIT=16'b1110111010111011;
    LogicCell40 value_cnt_11_LC_7_6_0 (
            .in0(N__2252),
            .in1(N__2275),
            .in2(_gnd_net_),
            .in3(N__2283),
            .lcout(value_cntZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2118),
            .ce(N__2085),
            .sr(N__2059));
    defparam value_cnt_9_LC_7_6_2.C_ON=1'b0;
    defparam value_cnt_9_LC_7_6_2.SEQ_MODE=4'b1011;
    defparam value_cnt_9_LC_7_6_2.LUT_INIT=16'b1111101010101111;
    LogicCell40 value_cnt_9_LC_7_6_2 (
            .in0(N__2253),
            .in1(_gnd_net_),
            .in2(N__2151),
            .in3(N__2140),
            .lcout(value_cntZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2118),
            .ce(N__2085),
            .sr(N__2059));
endmodule // incremental
