-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Mar 17 2018 18:15:53

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "incremental" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of incremental
entity incremental is
port (
    leds : out std_logic_vector(7 downto 0);
    reset : in std_logic;
    clk : in std_logic);
end incremental;

-- Architecture of incremental
-- View name is \INTERFACE\
architecture \INTERFACE\ of incremental is

signal \N__2704\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2674\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2665\ : std_logic;
signal \N__2664\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2655\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2638\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2619\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2550\ : std_logic;
signal \N__2547\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2526\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2524\ : std_logic;
signal \N__2523\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2521\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2505\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2502\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2491\ : std_logic;
signal \N__2490\ : std_logic;
signal \N__2487\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2467\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2448\ : std_logic;
signal \N__2447\ : std_logic;
signal \N__2446\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2438\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2424\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2417\ : std_logic;
signal \N__2416\ : std_logic;
signal \N__2413\ : std_logic;
signal \N__2408\ : std_logic;
signal \N__2403\ : std_logic;
signal \N__2400\ : std_logic;
signal \N__2397\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2379\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2377\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2373\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2351\ : std_logic;
signal \N__2350\ : std_logic;
signal \N__2349\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2346\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2343\ : std_logic;
signal \N__2342\ : std_logic;
signal \N__2341\ : std_logic;
signal \N__2340\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2338\ : std_logic;
signal \N__2337\ : std_logic;
signal \N__2336\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2321\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2305\ : std_logic;
signal \N__2296\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2277\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2275\ : std_logic;
signal \N__2272\ : std_logic;
signal \N__2269\ : std_logic;
signal \N__2266\ : std_logic;
signal \N__2263\ : std_logic;
signal \N__2260\ : std_logic;
signal \N__2253\ : std_logic;
signal \N__2252\ : std_logic;
signal \N__2247\ : std_logic;
signal \N__2246\ : std_logic;
signal \N__2245\ : std_logic;
signal \N__2244\ : std_logic;
signal \N__2243\ : std_logic;
signal \N__2242\ : std_logic;
signal \N__2241\ : std_logic;
signal \N__2240\ : std_logic;
signal \N__2239\ : std_logic;
signal \N__2238\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2236\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2233\ : std_logic;
signal \N__2230\ : std_logic;
signal \N__2215\ : std_logic;
signal \N__2214\ : std_logic;
signal \N__2199\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2197\ : std_logic;
signal \N__2196\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2194\ : std_logic;
signal \N__2193\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2189\ : std_logic;
signal \N__2186\ : std_logic;
signal \N__2183\ : std_logic;
signal \N__2180\ : std_logic;
signal \N__2175\ : std_logic;
signal \N__2164\ : std_logic;
signal \N__2151\ : std_logic;
signal \N__2148\ : std_logic;
signal \N__2145\ : std_logic;
signal \N__2142\ : std_logic;
signal \N__2141\ : std_logic;
signal \N__2140\ : std_logic;
signal \N__2137\ : std_logic;
signal \N__2134\ : std_logic;
signal \N__2131\ : std_logic;
signal \N__2128\ : std_logic;
signal \N__2125\ : std_logic;
signal \N__2118\ : std_logic;
signal \N__2117\ : std_logic;
signal \N__2116\ : std_logic;
signal \N__2115\ : std_logic;
signal \N__2114\ : std_logic;
signal \N__2113\ : std_logic;
signal \N__2112\ : std_logic;
signal \N__2111\ : std_logic;
signal \N__2110\ : std_logic;
signal \N__2091\ : std_logic;
signal \N__2088\ : std_logic;
signal \N__2085\ : std_logic;
signal \N__2084\ : std_logic;
signal \N__2083\ : std_logic;
signal \N__2082\ : std_logic;
signal \N__2081\ : std_logic;
signal \N__2070\ : std_logic;
signal \N__2067\ : std_logic;
signal \N__2064\ : std_logic;
signal \N__2063\ : std_logic;
signal \N__2062\ : std_logic;
signal \N__2061\ : std_logic;
signal \N__2060\ : std_logic;
signal \N__2059\ : std_logic;
signal \N__2058\ : std_logic;
signal \N__2057\ : std_logic;
signal \N__2056\ : std_logic;
signal \N__2037\ : std_logic;
signal \N__2034\ : std_logic;
signal \N__2031\ : std_logic;
signal \N__2030\ : std_logic;
signal \N__2027\ : std_logic;
signal \N__2026\ : std_logic;
signal \N__2023\ : std_logic;
signal \N__2020\ : std_logic;
signal \N__2017\ : std_logic;
signal \N__2010\ : std_logic;
signal \N__2007\ : std_logic;
signal \N__2004\ : std_logic;
signal \N__2001\ : std_logic;
signal \N__2000\ : std_logic;
signal \N__1999\ : std_logic;
signal \N__1996\ : std_logic;
signal \N__1993\ : std_logic;
signal \N__1990\ : std_logic;
signal \N__1983\ : std_logic;
signal \N__1980\ : std_logic;
signal \N__1977\ : std_logic;
signal \N__1974\ : std_logic;
signal \N__1971\ : std_logic;
signal \N__1970\ : std_logic;
signal \N__1967\ : std_logic;
signal \N__1964\ : std_logic;
signal \N__1961\ : std_logic;
signal \N__1956\ : std_logic;
signal \N__1953\ : std_logic;
signal \N__1950\ : std_logic;
signal \N__1947\ : std_logic;
signal \N__1946\ : std_logic;
signal \N__1945\ : std_logic;
signal \N__1942\ : std_logic;
signal \N__1937\ : std_logic;
signal \N__1932\ : std_logic;
signal \N__1929\ : std_logic;
signal \N__1928\ : std_logic;
signal \N__1927\ : std_logic;
signal \N__1922\ : std_logic;
signal \N__1919\ : std_logic;
signal \N__1914\ : std_logic;
signal \N__1911\ : std_logic;
signal \N__1908\ : std_logic;
signal \N__1907\ : std_logic;
signal \N__1906\ : std_logic;
signal \N__1903\ : std_logic;
signal \N__1900\ : std_logic;
signal \N__1897\ : std_logic;
signal \N__1890\ : std_logic;
signal \N__1887\ : std_logic;
signal \N__1884\ : std_logic;
signal \N__1881\ : std_logic;
signal \N__1880\ : std_logic;
signal \N__1879\ : std_logic;
signal \N__1876\ : std_logic;
signal \N__1873\ : std_logic;
signal \N__1870\ : std_logic;
signal \N__1863\ : std_logic;
signal \N__1862\ : std_logic;
signal \N__1861\ : std_logic;
signal \N__1858\ : std_logic;
signal \N__1855\ : std_logic;
signal \N__1852\ : std_logic;
signal \N__1849\ : std_logic;
signal \N__1842\ : std_logic;
signal \N__1839\ : std_logic;
signal \N__1836\ : std_logic;
signal \N__1833\ : std_logic;
signal \N__1832\ : std_logic;
signal \N__1831\ : std_logic;
signal \N__1828\ : std_logic;
signal \N__1825\ : std_logic;
signal \N__1822\ : std_logic;
signal \N__1819\ : std_logic;
signal \N__1816\ : std_logic;
signal \N__1809\ : std_logic;
signal \N__1806\ : std_logic;
signal \N__1803\ : std_logic;
signal \N__1800\ : std_logic;
signal \N__1799\ : std_logic;
signal \N__1798\ : std_logic;
signal \N__1795\ : std_logic;
signal \N__1792\ : std_logic;
signal \N__1789\ : std_logic;
signal \N__1786\ : std_logic;
signal \N__1779\ : std_logic;
signal \N__1776\ : std_logic;
signal \N__1773\ : std_logic;
signal \N__1770\ : std_logic;
signal \N__1769\ : std_logic;
signal \N__1768\ : std_logic;
signal \N__1765\ : std_logic;
signal \N__1762\ : std_logic;
signal \N__1759\ : std_logic;
signal \N__1756\ : std_logic;
signal \N__1749\ : std_logic;
signal \N__1746\ : std_logic;
signal \N__1743\ : std_logic;
signal \N__1740\ : std_logic;
signal \N__1739\ : std_logic;
signal \N__1736\ : std_logic;
signal \N__1735\ : std_logic;
signal \N__1732\ : std_logic;
signal \N__1729\ : std_logic;
signal \N__1726\ : std_logic;
signal \N__1719\ : std_logic;
signal \N__1716\ : std_logic;
signal \N__1713\ : std_logic;
signal \N__1710\ : std_logic;
signal \N__1709\ : std_logic;
signal \N__1708\ : std_logic;
signal \N__1705\ : std_logic;
signal \N__1702\ : std_logic;
signal \N__1699\ : std_logic;
signal \N__1696\ : std_logic;
signal \N__1693\ : std_logic;
signal \N__1686\ : std_logic;
signal \N__1683\ : std_logic;
signal \N__1680\ : std_logic;
signal \N__1677\ : std_logic;
signal \N__1676\ : std_logic;
signal \N__1673\ : std_logic;
signal \N__1672\ : std_logic;
signal \N__1669\ : std_logic;
signal \N__1666\ : std_logic;
signal \N__1663\ : std_logic;
signal \N__1656\ : std_logic;
signal \N__1653\ : std_logic;
signal \N__1650\ : std_logic;
signal \N__1647\ : std_logic;
signal \N__1646\ : std_logic;
signal \N__1645\ : std_logic;
signal \N__1642\ : std_logic;
signal \N__1639\ : std_logic;
signal \N__1636\ : std_logic;
signal \N__1633\ : std_logic;
signal \N__1626\ : std_logic;
signal \N__1623\ : std_logic;
signal \N__1620\ : std_logic;
signal \N__1617\ : std_logic;
signal \N__1616\ : std_logic;
signal \N__1615\ : std_logic;
signal \N__1612\ : std_logic;
signal \N__1609\ : std_logic;
signal \N__1606\ : std_logic;
signal \N__1603\ : std_logic;
signal \N__1596\ : std_logic;
signal \N__1593\ : std_logic;
signal \N__1590\ : std_logic;
signal \N__1587\ : std_logic;
signal \N__1586\ : std_logic;
signal \N__1585\ : std_logic;
signal \N__1582\ : std_logic;
signal \N__1579\ : std_logic;
signal \N__1576\ : std_logic;
signal \N__1573\ : std_logic;
signal \N__1570\ : std_logic;
signal \N__1563\ : std_logic;
signal \N__1560\ : std_logic;
signal \N__1557\ : std_logic;
signal \N__1554\ : std_logic;
signal \N__1553\ : std_logic;
signal \N__1552\ : std_logic;
signal \N__1549\ : std_logic;
signal \N__1546\ : std_logic;
signal \N__1543\ : std_logic;
signal \N__1540\ : std_logic;
signal \N__1533\ : std_logic;
signal \N__1530\ : std_logic;
signal \N__1527\ : std_logic;
signal \N__1524\ : std_logic;
signal \N__1523\ : std_logic;
signal \N__1522\ : std_logic;
signal \N__1519\ : std_logic;
signal \N__1516\ : std_logic;
signal \N__1513\ : std_logic;
signal \N__1510\ : std_logic;
signal \N__1503\ : std_logic;
signal \N__1500\ : std_logic;
signal \N__1497\ : std_logic;
signal \N__1494\ : std_logic;
signal \N__1491\ : std_logic;
signal \N__1490\ : std_logic;
signal \N__1489\ : std_logic;
signal \N__1486\ : std_logic;
signal \N__1483\ : std_logic;
signal \N__1480\ : std_logic;
signal \N__1477\ : std_logic;
signal \N__1474\ : std_logic;
signal \N__1467\ : std_logic;
signal \N__1464\ : std_logic;
signal \N__1461\ : std_logic;
signal \N__1458\ : std_logic;
signal \N__1455\ : std_logic;
signal \N__1454\ : std_logic;
signal \N__1453\ : std_logic;
signal \N__1450\ : std_logic;
signal \N__1447\ : std_logic;
signal \N__1444\ : std_logic;
signal \N__1441\ : std_logic;
signal \N__1434\ : std_logic;
signal \N__1431\ : std_logic;
signal \N__1428\ : std_logic;
signal \N__1425\ : std_logic;
signal \N__1424\ : std_logic;
signal \N__1419\ : std_logic;
signal \N__1416\ : std_logic;
signal \N__1413\ : std_logic;
signal \N__1410\ : std_logic;
signal \N__1409\ : std_logic;
signal \N__1404\ : std_logic;
signal \N__1401\ : std_logic;
signal \N__1400\ : std_logic;
signal \N__1399\ : std_logic;
signal \N__1396\ : std_logic;
signal \N__1393\ : std_logic;
signal \N__1390\ : std_logic;
signal \N__1383\ : std_logic;
signal \N__1382\ : std_logic;
signal \N__1381\ : std_logic;
signal \N__1378\ : std_logic;
signal \N__1375\ : std_logic;
signal \N__1372\ : std_logic;
signal \N__1365\ : std_logic;
signal \N__1364\ : std_logic;
signal \N__1363\ : std_logic;
signal \N__1360\ : std_logic;
signal \N__1357\ : std_logic;
signal \N__1354\ : std_logic;
signal \N__1351\ : std_logic;
signal \N__1344\ : std_logic;
signal \N__1341\ : std_logic;
signal \N__1338\ : std_logic;
signal \N__1335\ : std_logic;
signal \N__1334\ : std_logic;
signal \N__1333\ : std_logic;
signal \N__1330\ : std_logic;
signal \N__1327\ : std_logic;
signal \N__1324\ : std_logic;
signal \N__1321\ : std_logic;
signal \N__1318\ : std_logic;
signal \N__1311\ : std_logic;
signal \N__1308\ : std_logic;
signal \N__1305\ : std_logic;
signal \N__1302\ : std_logic;
signal \N__1301\ : std_logic;
signal \N__1300\ : std_logic;
signal \N__1297\ : std_logic;
signal \N__1294\ : std_logic;
signal \N__1291\ : std_logic;
signal \N__1288\ : std_logic;
signal \N__1281\ : std_logic;
signal \N__1278\ : std_logic;
signal \N__1275\ : std_logic;
signal \N__1272\ : std_logic;
signal \N__1271\ : std_logic;
signal \N__1270\ : std_logic;
signal \N__1267\ : std_logic;
signal \N__1264\ : std_logic;
signal \N__1261\ : std_logic;
signal \N__1258\ : std_logic;
signal \N__1251\ : std_logic;
signal \N__1248\ : std_logic;
signal \N__1245\ : std_logic;
signal \N__1242\ : std_logic;
signal \N__1241\ : std_logic;
signal \N__1240\ : std_logic;
signal \N__1237\ : std_logic;
signal \N__1234\ : std_logic;
signal \N__1231\ : std_logic;
signal \N__1224\ : std_logic;
signal \N__1223\ : std_logic;
signal \N__1220\ : std_logic;
signal \N__1217\ : std_logic;
signal \N__1212\ : std_logic;
signal \N__1211\ : std_logic;
signal \N__1210\ : std_logic;
signal \N__1207\ : std_logic;
signal \N__1204\ : std_logic;
signal \N__1203\ : std_logic;
signal \N__1194\ : std_logic;
signal \N__1191\ : std_logic;
signal \N__1190\ : std_logic;
signal \N__1189\ : std_logic;
signal \N__1186\ : std_logic;
signal \N__1185\ : std_logic;
signal \N__1180\ : std_logic;
signal \N__1175\ : std_logic;
signal \N__1170\ : std_logic;
signal \N__1169\ : std_logic;
signal \N__1168\ : std_logic;
signal \N__1163\ : std_logic;
signal \N__1160\ : std_logic;
signal \N__1155\ : std_logic;
signal \N__1154\ : std_logic;
signal \N__1153\ : std_logic;
signal \N__1150\ : std_logic;
signal \N__1145\ : std_logic;
signal \N__1142\ : std_logic;
signal \N__1137\ : std_logic;
signal \N__1134\ : std_logic;
signal \N__1131\ : std_logic;
signal \N__1128\ : std_logic;
signal \N__1125\ : std_logic;
signal \N__1122\ : std_logic;
signal \N__1119\ : std_logic;
signal \N__1116\ : std_logic;
signal \N__1113\ : std_logic;
signal \N__1110\ : std_logic;
signal \N__1107\ : std_logic;
signal \N__1104\ : std_logic;
signal \N__1101\ : std_logic;
signal \N__1098\ : std_logic;
signal \N__1095\ : std_logic;
signal \N__1092\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \op_eq_un4_fin_cnt_20_3_cascade_\ : std_logic;
signal op_eq_un4_fin_cnt_20_4 : std_logic;
signal op_eq_un4_fin_cnt_21_9 : std_logic;
signal op_eq_un4_fin_cnt_21_11 : std_logic;
signal op_eq_un4_fin_cnt_21_10 : std_logic;
signal op_eq_un4_fin_cnt_21_8 : std_logic;
signal op_eq_un4_fin_cnt_20 : std_logic;
signal op_eq_un4_fin_cnt_21 : std_logic;
signal \UC.epZ0Z_3\ : std_logic;
signal \UC.epZ0Z_6\ : std_logic;
signal \UC.value_cnte_0_i\ : std_logic;
signal \UC.epZ0Z_4\ : std_logic;
signal \UC.sr_reg\ : std_logic;
signal \UC.epZ0Z_0\ : std_logic;
signal \UC.epZ0Z_8\ : std_logic;
signal \UC.epZ0Z_1\ : std_logic;
signal \UC.epZ0Z_7\ : std_logic;
signal \value_cntZ0Z_0\ : std_logic;
signal \bfn_6_5_0_\ : std_logic;
signal \value_cntZ0Z_1\ : std_logic;
signal \value_cnt_cry_0_THRU_CO\ : std_logic;
signal value_cnt_cry_0 : std_logic;
signal \value_cntZ0Z_2\ : std_logic;
signal \value_cnt_cry_1_THRU_CO\ : std_logic;
signal value_cnt_cry_1 : std_logic;
signal \value_cntZ0Z_3\ : std_logic;
signal \value_cnt_cry_2_THRU_CO\ : std_logic;
signal value_cnt_cry_2 : std_logic;
signal \value_cntZ0Z_4\ : std_logic;
signal \value_cnt_cry_3_THRU_CO\ : std_logic;
signal value_cnt_cry_3 : std_logic;
signal \value_cntZ0Z_5\ : std_logic;
signal \value_cnt_cry_4_THRU_CO\ : std_logic;
signal value_cnt_cry_4 : std_logic;
signal \value_cntZ0Z_6\ : std_logic;
signal \value_cnt_cry_5_THRU_CO\ : std_logic;
signal value_cnt_cry_5 : std_logic;
signal \value_cntZ0Z_7\ : std_logic;
signal \value_cnt_cry_6_THRU_CO\ : std_logic;
signal value_cnt_cry_6 : std_logic;
signal value_cnt_cry_7 : std_logic;
signal \value_cntZ0Z_8\ : std_logic;
signal \value_cnt_cry_7_THRU_CO\ : std_logic;
signal \bfn_6_6_0_\ : std_logic;
signal value_cnt_cry_8 : std_logic;
signal \value_cntZ0Z_10\ : std_logic;
signal \value_cnt_cry_9_THRU_CO\ : std_logic;
signal value_cnt_cry_9 : std_logic;
signal value_cnt_cry_10 : std_logic;
signal \value_cntZ0Z_12\ : std_logic;
signal \value_cnt_cry_11_THRU_CO\ : std_logic;
signal value_cnt_cry_11 : std_logic;
signal \value_cntZ0Z_13\ : std_logic;
signal \value_cnt_cry_12_THRU_CO\ : std_logic;
signal value_cnt_cry_12 : std_logic;
signal \value_cntZ0Z_14\ : std_logic;
signal \value_cnt_cry_13_THRU_CO\ : std_logic;
signal value_cnt_cry_13 : std_logic;
signal \value_cntZ0Z_15\ : std_logic;
signal \value_cnt_cry_14_THRU_CO\ : std_logic;
signal value_cnt_cry_14 : std_logic;
signal value_cnt_cry_15 : std_logic;
signal \value_cntZ0Z_16\ : std_logic;
signal \value_cnt_cry_15_THRU_CO\ : std_logic;
signal \bfn_6_7_0_\ : std_logic;
signal \value_cntZ0Z_17\ : std_logic;
signal \value_cnt_cry_16_THRU_CO\ : std_logic;
signal value_cnt_cry_16 : std_logic;
signal \value_cntZ0Z_18\ : std_logic;
signal \value_cnt_cry_17_THRU_CO\ : std_logic;
signal value_cnt_cry_17 : std_logic;
signal \value_cntZ0Z_19\ : std_logic;
signal \value_cnt_cry_18_THRU_CO\ : std_logic;
signal value_cnt_cry_18 : std_logic;
signal \value_cntZ0Z_20\ : std_logic;
signal \value_cnt_cry_19_THRU_CO\ : std_logic;
signal value_cnt_cry_19 : std_logic;
signal \value_cntZ0Z_21\ : std_logic;
signal \value_cnt_cry_20_THRU_CO\ : std_logic;
signal value_cnt_cry_20 : std_logic;
signal \value_cntZ0Z_22\ : std_logic;
signal \value_cnt_cry_21_THRU_CO\ : std_logic;
signal value_cnt_cry_21 : std_logic;
signal value_cnt_cry_22 : std_logic;
signal \value_cntZ0Z_23\ : std_logic;
signal leds_c_0 : std_logic;
signal \register10Z0Z_0\ : std_logic;
signal leds_c_1 : std_logic;
signal leds_c_2 : std_logic;
signal leds_c_3 : std_logic;
signal leds_c_4 : std_logic;
signal leds_c_5 : std_logic;
signal sl_reg : std_logic;
signal \register10Z0Z_9\ : std_logic;
signal leds_c_6 : std_logic;
signal leds_c_7 : std_logic;
signal un1_sr_reg_0_i : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \value_cnt_cry_10_THRU_CO\ : std_logic;
signal \value_cntZ0Z_11\ : std_logic;
signal \UC_un1_ld_cnt_0_i\ : std_logic;
signal \value_cnt_cry_8_THRU_CO\ : std_logic;
signal \value_cntZ0Z_9\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_c_g : std_logic;
signal value_cnte_0_i_g : std_logic;
signal reset_c_g : std_logic;

signal reset_wire : std_logic;
signal clk_wire : std_logic;
signal leds_wire : std_logic_vector(7 downto 0);

begin
    reset_wire <= reset;
    clk_wire <= clk;
    leds <= leds_wire;

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__2702\,
            GLOBALBUFFEROUTPUT => reset_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2704\,
            DIN => \N__2703\,
            DOUT => \N__2702\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2704\,
            PADOUT => \N__2703\,
            PADIN => \N__2702\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__2692\,
            GLOBALBUFFEROUTPUT => clk_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2694\,
            DIN => \N__2693\,
            DOUT => \N__2692\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2694\,
            PADOUT => \N__2693\,
            PADIN => \N__2692\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2683\,
            DIN => \N__2682\,
            DOUT => \N__2681\,
            PACKAGEPIN => leds_wire(1)
        );

    \leds_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2683\,
            PADOUT => \N__2682\,
            PADIN => \N__2681\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1914\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2674\,
            DIN => \N__2673\,
            DOUT => \N__2672\,
            PACKAGEPIN => leds_wire(5)
        );

    \leds_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2674\,
            PADOUT => \N__2673\,
            PADIN => \N__2672\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2550\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2665\,
            DIN => \N__2664\,
            DOUT => \N__2663\,
            PACKAGEPIN => leds_wire(0)
        );

    \leds_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2665\,
            PADOUT => \N__2664\,
            PADIN => \N__2663\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1956\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2656\,
            DIN => \N__2655\,
            DOUT => \N__2654\,
            PACKAGEPIN => leds_wire(4)
        );

    \leds_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2656\,
            PADOUT => \N__2655\,
            PADIN => \N__2654\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2574\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2647\,
            DIN => \N__2646\,
            DOUT => \N__2645\,
            PACKAGEPIN => leds_wire(3)
        );

    \leds_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2647\,
            PADOUT => \N__2646\,
            PADIN => \N__2645\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2601\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2638\,
            DIN => \N__2637\,
            DOUT => \N__2636\,
            PACKAGEPIN => leds_wire(7)
        );

    \leds_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2638\,
            PADOUT => \N__2637\,
            PADIN => \N__2636\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2433\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2629\,
            DIN => \N__2628\,
            DOUT => \N__2627\,
            PACKAGEPIN => leds_wire(2)
        );

    \leds_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2629\,
            PADOUT => \N__2628\,
            PADIN => \N__2627\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1890\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \leds_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2620\,
            DIN => \N__2619\,
            DOUT => \N__2618\,
            PACKAGEPIN => leds_wire(6)
        );

    \leds_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2620\,
            PADOUT => \N__2619\,
            PADIN => \N__2618\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2454\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__598\ : IoInMux
    port map (
            O => \N__2601\,
            I => \N__2598\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__2598\,
            I => \N__2595\
        );

    \I__596\ : IoSpan4Mux
    port map (
            O => \N__2595\,
            I => \N__2591\
        );

    \I__595\ : CascadeMux
    port map (
            O => \N__2594\,
            I => \N__2588\
        );

    \I__594\ : Span4Mux_s3_h
    port map (
            O => \N__2591\,
            I => \N__2584\
        );

    \I__593\ : InMux
    port map (
            O => \N__2588\,
            I => \N__2579\
        );

    \I__592\ : InMux
    port map (
            O => \N__2587\,
            I => \N__2579\
        );

    \I__591\ : Odrv4
    port map (
            O => \N__2584\,
            I => leds_c_3
        );

    \I__590\ : LocalMux
    port map (
            O => \N__2579\,
            I => leds_c_3
        );

    \I__589\ : IoInMux
    port map (
            O => \N__2574\,
            I => \N__2571\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__2571\,
            I => \N__2567\
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__2570\,
            I => \N__2564\
        );

    \I__586\ : Span12Mux_s6_h
    port map (
            O => \N__2567\,
            I => \N__2560\
        );

    \I__585\ : InMux
    port map (
            O => \N__2564\,
            I => \N__2555\
        );

    \I__584\ : InMux
    port map (
            O => \N__2563\,
            I => \N__2555\
        );

    \I__583\ : Odrv12
    port map (
            O => \N__2560\,
            I => leds_c_4
        );

    \I__582\ : LocalMux
    port map (
            O => \N__2555\,
            I => leds_c_4
        );

    \I__581\ : IoInMux
    port map (
            O => \N__2550\,
            I => \N__2547\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__2547\,
            I => \N__2544\
        );

    \I__579\ : Span4Mux_s3_h
    port map (
            O => \N__2544\,
            I => \N__2541\
        );

    \I__578\ : Span4Mux_v
    port map (
            O => \N__2541\,
            I => \N__2536\
        );

    \I__577\ : InMux
    port map (
            O => \N__2540\,
            I => \N__2531\
        );

    \I__576\ : InMux
    port map (
            O => \N__2539\,
            I => \N__2531\
        );

    \I__575\ : Odrv4
    port map (
            O => \N__2536\,
            I => leds_c_5
        );

    \I__574\ : LocalMux
    port map (
            O => \N__2531\,
            I => leds_c_5
        );

    \I__573\ : InMux
    port map (
            O => \N__2526\,
            I => \N__2505\
        );

    \I__572\ : InMux
    port map (
            O => \N__2525\,
            I => \N__2505\
        );

    \I__571\ : InMux
    port map (
            O => \N__2524\,
            I => \N__2505\
        );

    \I__570\ : InMux
    port map (
            O => \N__2523\,
            I => \N__2505\
        );

    \I__569\ : InMux
    port map (
            O => \N__2522\,
            I => \N__2505\
        );

    \I__568\ : InMux
    port map (
            O => \N__2521\,
            I => \N__2505\
        );

    \I__567\ : InMux
    port map (
            O => \N__2520\,
            I => \N__2505\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__2505\,
            I => \N__2498\
        );

    \I__565\ : InMux
    port map (
            O => \N__2504\,
            I => \N__2491\
        );

    \I__564\ : InMux
    port map (
            O => \N__2503\,
            I => \N__2491\
        );

    \I__563\ : InMux
    port map (
            O => \N__2502\,
            I => \N__2491\
        );

    \I__562\ : InMux
    port map (
            O => \N__2501\,
            I => \N__2487\
        );

    \I__561\ : Span4Mux_v
    port map (
            O => \N__2498\,
            I => \N__2484\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__2491\,
            I => \N__2481\
        );

    \I__559\ : InMux
    port map (
            O => \N__2490\,
            I => \N__2478\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__2487\,
            I => sl_reg
        );

    \I__557\ : Odrv4
    port map (
            O => \N__2484\,
            I => sl_reg
        );

    \I__556\ : Odrv4
    port map (
            O => \N__2481\,
            I => sl_reg
        );

    \I__555\ : LocalMux
    port map (
            O => \N__2478\,
            I => sl_reg
        );

    \I__554\ : InMux
    port map (
            O => \N__2469\,
            I => \N__2462\
        );

    \I__553\ : InMux
    port map (
            O => \N__2468\,
            I => \N__2462\
        );

    \I__552\ : InMux
    port map (
            O => \N__2467\,
            I => \N__2459\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__2462\,
            I => \register10Z0Z_9\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__2459\,
            I => \register10Z0Z_9\
        );

    \I__549\ : IoInMux
    port map (
            O => \N__2454\,
            I => \N__2451\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__2451\,
            I => \N__2448\
        );

    \I__547\ : Span12Mux_s6_h
    port map (
            O => \N__2448\,
            I => \N__2443\
        );

    \I__546\ : InMux
    port map (
            O => \N__2447\,
            I => \N__2438\
        );

    \I__545\ : InMux
    port map (
            O => \N__2446\,
            I => \N__2438\
        );

    \I__544\ : Odrv12
    port map (
            O => \N__2443\,
            I => leds_c_6
        );

    \I__543\ : LocalMux
    port map (
            O => \N__2438\,
            I => leds_c_6
        );

    \I__542\ : IoInMux
    port map (
            O => \N__2433\,
            I => \N__2430\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__2430\,
            I => \N__2427\
        );

    \I__540\ : IoSpan4Mux
    port map (
            O => \N__2427\,
            I => \N__2424\
        );

    \I__539\ : Span4Mux_s3_h
    port map (
            O => \N__2424\,
            I => \N__2420\
        );

    \I__538\ : CascadeMux
    port map (
            O => \N__2423\,
            I => \N__2417\
        );

    \I__537\ : Span4Mux_v
    port map (
            O => \N__2420\,
            I => \N__2413\
        );

    \I__536\ : InMux
    port map (
            O => \N__2417\,
            I => \N__2408\
        );

    \I__535\ : InMux
    port map (
            O => \N__2416\,
            I => \N__2408\
        );

    \I__534\ : Odrv4
    port map (
            O => \N__2413\,
            I => leds_c_7
        );

    \I__533\ : LocalMux
    port map (
            O => \N__2408\,
            I => leds_c_7
        );

    \I__532\ : CEMux
    port map (
            O => \N__2403\,
            I => \N__2400\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__2400\,
            I => \N__2397\
        );

    \I__530\ : Span4Mux_v
    port map (
            O => \N__2397\,
            I => \N__2393\
        );

    \I__529\ : CEMux
    port map (
            O => \N__2396\,
            I => \N__2390\
        );

    \I__528\ : Span4Mux_h
    port map (
            O => \N__2393\,
            I => \N__2387\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__2390\,
            I => \N__2384\
        );

    \I__526\ : Odrv4
    port map (
            O => \N__2387\,
            I => un1_sr_reg_0_i
        );

    \I__525\ : Odrv12
    port map (
            O => \N__2384\,
            I => un1_sr_reg_0_i
        );

    \I__524\ : CascadeMux
    port map (
            O => \N__2379\,
            I => \N__2373\
        );

    \I__523\ : InMux
    port map (
            O => \N__2378\,
            I => \N__2363\
        );

    \I__522\ : InMux
    port map (
            O => \N__2377\,
            I => \N__2363\
        );

    \I__521\ : InMux
    port map (
            O => \N__2376\,
            I => \N__2363\
        );

    \I__520\ : InMux
    port map (
            O => \N__2373\,
            I => \N__2354\
        );

    \I__519\ : InMux
    port map (
            O => \N__2372\,
            I => \N__2354\
        );

    \I__518\ : InMux
    port map (
            O => \N__2371\,
            I => \N__2354\
        );

    \I__517\ : InMux
    port map (
            O => \N__2370\,
            I => \N__2354\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__2363\,
            I => \N__2351\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__2354\,
            I => \N__2333\
        );

    \I__514\ : Span4Mux_v
    port map (
            O => \N__2351\,
            I => \N__2330\
        );

    \I__513\ : InMux
    port map (
            O => \N__2350\,
            I => \N__2321\
        );

    \I__512\ : InMux
    port map (
            O => \N__2349\,
            I => \N__2321\
        );

    \I__511\ : InMux
    port map (
            O => \N__2348\,
            I => \N__2321\
        );

    \I__510\ : InMux
    port map (
            O => \N__2347\,
            I => \N__2321\
        );

    \I__509\ : InMux
    port map (
            O => \N__2346\,
            I => \N__2312\
        );

    \I__508\ : InMux
    port map (
            O => \N__2345\,
            I => \N__2312\
        );

    \I__507\ : InMux
    port map (
            O => \N__2344\,
            I => \N__2312\
        );

    \I__506\ : InMux
    port map (
            O => \N__2343\,
            I => \N__2312\
        );

    \I__505\ : InMux
    port map (
            O => \N__2342\,
            I => \N__2305\
        );

    \I__504\ : InMux
    port map (
            O => \N__2341\,
            I => \N__2305\
        );

    \I__503\ : InMux
    port map (
            O => \N__2340\,
            I => \N__2305\
        );

    \I__502\ : InMux
    port map (
            O => \N__2339\,
            I => \N__2296\
        );

    \I__501\ : InMux
    port map (
            O => \N__2338\,
            I => \N__2296\
        );

    \I__500\ : InMux
    port map (
            O => \N__2337\,
            I => \N__2296\
        );

    \I__499\ : InMux
    port map (
            O => \N__2336\,
            I => \N__2296\
        );

    \I__498\ : Odrv4
    port map (
            O => \N__2333\,
            I => \CONSTANT_ONE_NET\
        );

    \I__497\ : Odrv4
    port map (
            O => \N__2330\,
            I => \CONSTANT_ONE_NET\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__2321\,
            I => \CONSTANT_ONE_NET\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__2312\,
            I => \CONSTANT_ONE_NET\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__2305\,
            I => \CONSTANT_ONE_NET\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__2296\,
            I => \CONSTANT_ONE_NET\
        );

    \I__492\ : InMux
    port map (
            O => \N__2283\,
            I => \N__2280\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__2280\,
            I => \value_cnt_cry_10_THRU_CO\
        );

    \I__490\ : InMux
    port map (
            O => \N__2277\,
            I => \N__2272\
        );

    \I__489\ : CascadeMux
    port map (
            O => \N__2276\,
            I => \N__2269\
        );

    \I__488\ : InMux
    port map (
            O => \N__2275\,
            I => \N__2266\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__2272\,
            I => \N__2263\
        );

    \I__486\ : InMux
    port map (
            O => \N__2269\,
            I => \N__2260\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__2266\,
            I => \value_cntZ0Z_11\
        );

    \I__484\ : Odrv12
    port map (
            O => \N__2263\,
            I => \value_cntZ0Z_11\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__2260\,
            I => \value_cntZ0Z_11\
        );

    \I__482\ : InMux
    port map (
            O => \N__2253\,
            I => \N__2247\
        );

    \I__481\ : InMux
    port map (
            O => \N__2252\,
            I => \N__2247\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__2247\,
            I => \N__2230\
        );

    \I__479\ : InMux
    port map (
            O => \N__2246\,
            I => \N__2215\
        );

    \I__478\ : InMux
    port map (
            O => \N__2245\,
            I => \N__2215\
        );

    \I__477\ : InMux
    port map (
            O => \N__2244\,
            I => \N__2215\
        );

    \I__476\ : InMux
    port map (
            O => \N__2243\,
            I => \N__2215\
        );

    \I__475\ : InMux
    port map (
            O => \N__2242\,
            I => \N__2215\
        );

    \I__474\ : InMux
    port map (
            O => \N__2241\,
            I => \N__2215\
        );

    \I__473\ : InMux
    port map (
            O => \N__2240\,
            I => \N__2215\
        );

    \I__472\ : InMux
    port map (
            O => \N__2239\,
            I => \N__2199\
        );

    \I__471\ : InMux
    port map (
            O => \N__2238\,
            I => \N__2199\
        );

    \I__470\ : InMux
    port map (
            O => \N__2237\,
            I => \N__2199\
        );

    \I__469\ : InMux
    port map (
            O => \N__2236\,
            I => \N__2199\
        );

    \I__468\ : InMux
    port map (
            O => \N__2235\,
            I => \N__2199\
        );

    \I__467\ : InMux
    port map (
            O => \N__2234\,
            I => \N__2199\
        );

    \I__466\ : InMux
    port map (
            O => \N__2233\,
            I => \N__2199\
        );

    \I__465\ : Span4Mux_h
    port map (
            O => \N__2230\,
            I => \N__2189\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__2215\,
            I => \N__2186\
        );

    \I__463\ : InMux
    port map (
            O => \N__2214\,
            I => \N__2183\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__2199\,
            I => \N__2180\
        );

    \I__461\ : InMux
    port map (
            O => \N__2198\,
            I => \N__2175\
        );

    \I__460\ : InMux
    port map (
            O => \N__2197\,
            I => \N__2175\
        );

    \I__459\ : InMux
    port map (
            O => \N__2196\,
            I => \N__2164\
        );

    \I__458\ : InMux
    port map (
            O => \N__2195\,
            I => \N__2164\
        );

    \I__457\ : InMux
    port map (
            O => \N__2194\,
            I => \N__2164\
        );

    \I__456\ : InMux
    port map (
            O => \N__2193\,
            I => \N__2164\
        );

    \I__455\ : InMux
    port map (
            O => \N__2192\,
            I => \N__2164\
        );

    \I__454\ : Odrv4
    port map (
            O => \N__2189\,
            I => \UC_un1_ld_cnt_0_i\
        );

    \I__453\ : Odrv4
    port map (
            O => \N__2186\,
            I => \UC_un1_ld_cnt_0_i\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__2183\,
            I => \UC_un1_ld_cnt_0_i\
        );

    \I__451\ : Odrv4
    port map (
            O => \N__2180\,
            I => \UC_un1_ld_cnt_0_i\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__2175\,
            I => \UC_un1_ld_cnt_0_i\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2164\,
            I => \UC_un1_ld_cnt_0_i\
        );

    \I__448\ : CascadeMux
    port map (
            O => \N__2151\,
            I => \N__2148\
        );

    \I__447\ : InMux
    port map (
            O => \N__2148\,
            I => \N__2145\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__2145\,
            I => \value_cnt_cry_8_THRU_CO\
        );

    \I__445\ : InMux
    port map (
            O => \N__2142\,
            I => \N__2137\
        );

    \I__444\ : CascadeMux
    port map (
            O => \N__2141\,
            I => \N__2134\
        );

    \I__443\ : InMux
    port map (
            O => \N__2140\,
            I => \N__2131\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__2137\,
            I => \N__2128\
        );

    \I__441\ : InMux
    port map (
            O => \N__2134\,
            I => \N__2125\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__2131\,
            I => \value_cntZ0Z_9\
        );

    \I__439\ : Odrv12
    port map (
            O => \N__2128\,
            I => \value_cntZ0Z_9\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2125\,
            I => \value_cntZ0Z_9\
        );

    \I__437\ : ClkMux
    port map (
            O => \N__2118\,
            I => \N__2091\
        );

    \I__436\ : ClkMux
    port map (
            O => \N__2117\,
            I => \N__2091\
        );

    \I__435\ : ClkMux
    port map (
            O => \N__2116\,
            I => \N__2091\
        );

    \I__434\ : ClkMux
    port map (
            O => \N__2115\,
            I => \N__2091\
        );

    \I__433\ : ClkMux
    port map (
            O => \N__2114\,
            I => \N__2091\
        );

    \I__432\ : ClkMux
    port map (
            O => \N__2113\,
            I => \N__2091\
        );

    \I__431\ : ClkMux
    port map (
            O => \N__2112\,
            I => \N__2091\
        );

    \I__430\ : ClkMux
    port map (
            O => \N__2111\,
            I => \N__2091\
        );

    \I__429\ : ClkMux
    port map (
            O => \N__2110\,
            I => \N__2091\
        );

    \I__428\ : GlobalMux
    port map (
            O => \N__2091\,
            I => \N__2088\
        );

    \I__427\ : gio2CtrlBuf
    port map (
            O => \N__2088\,
            I => clk_c_g
        );

    \I__426\ : CEMux
    port map (
            O => \N__2085\,
            I => \N__2070\
        );

    \I__425\ : CEMux
    port map (
            O => \N__2084\,
            I => \N__2070\
        );

    \I__424\ : CEMux
    port map (
            O => \N__2083\,
            I => \N__2070\
        );

    \I__423\ : CEMux
    port map (
            O => \N__2082\,
            I => \N__2070\
        );

    \I__422\ : CEMux
    port map (
            O => \N__2081\,
            I => \N__2070\
        );

    \I__421\ : GlobalMux
    port map (
            O => \N__2070\,
            I => \N__2067\
        );

    \I__420\ : gio2CtrlBuf
    port map (
            O => \N__2067\,
            I => value_cnte_0_i_g
        );

    \I__419\ : SRMux
    port map (
            O => \N__2064\,
            I => \N__2037\
        );

    \I__418\ : SRMux
    port map (
            O => \N__2063\,
            I => \N__2037\
        );

    \I__417\ : SRMux
    port map (
            O => \N__2062\,
            I => \N__2037\
        );

    \I__416\ : SRMux
    port map (
            O => \N__2061\,
            I => \N__2037\
        );

    \I__415\ : SRMux
    port map (
            O => \N__2060\,
            I => \N__2037\
        );

    \I__414\ : SRMux
    port map (
            O => \N__2059\,
            I => \N__2037\
        );

    \I__413\ : SRMux
    port map (
            O => \N__2058\,
            I => \N__2037\
        );

    \I__412\ : SRMux
    port map (
            O => \N__2057\,
            I => \N__2037\
        );

    \I__411\ : SRMux
    port map (
            O => \N__2056\,
            I => \N__2037\
        );

    \I__410\ : GlobalMux
    port map (
            O => \N__2037\,
            I => \N__2034\
        );

    \I__409\ : gio2CtrlBuf
    port map (
            O => \N__2034\,
            I => reset_c_g
        );

    \I__408\ : CascadeMux
    port map (
            O => \N__2031\,
            I => \N__2027\
        );

    \I__407\ : InMux
    port map (
            O => \N__2030\,
            I => \N__2023\
        );

    \I__406\ : InMux
    port map (
            O => \N__2027\,
            I => \N__2020\
        );

    \I__405\ : InMux
    port map (
            O => \N__2026\,
            I => \N__2017\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__2023\,
            I => \value_cntZ0Z_21\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2020\,
            I => \value_cntZ0Z_21\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2017\,
            I => \value_cntZ0Z_21\
        );

    \I__401\ : InMux
    port map (
            O => \N__2010\,
            I => \N__2007\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__2007\,
            I => \value_cnt_cry_20_THRU_CO\
        );

    \I__399\ : InMux
    port map (
            O => \N__2004\,
            I => value_cnt_cry_20
        );

    \I__398\ : InMux
    port map (
            O => \N__2001\,
            I => \N__1996\
        );

    \I__397\ : InMux
    port map (
            O => \N__2000\,
            I => \N__1993\
        );

    \I__396\ : InMux
    port map (
            O => \N__1999\,
            I => \N__1990\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__1996\,
            I => \value_cntZ0Z_22\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__1993\,
            I => \value_cntZ0Z_22\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__1990\,
            I => \value_cntZ0Z_22\
        );

    \I__392\ : InMux
    port map (
            O => \N__1983\,
            I => \N__1980\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__1980\,
            I => \value_cnt_cry_21_THRU_CO\
        );

    \I__390\ : InMux
    port map (
            O => \N__1977\,
            I => value_cnt_cry_21
        );

    \I__389\ : InMux
    port map (
            O => \N__1974\,
            I => value_cnt_cry_22
        );

    \I__388\ : InMux
    port map (
            O => \N__1971\,
            I => \N__1967\
        );

    \I__387\ : InMux
    port map (
            O => \N__1970\,
            I => \N__1964\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__1967\,
            I => \N__1961\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__1964\,
            I => \value_cntZ0Z_23\
        );

    \I__384\ : Odrv4
    port map (
            O => \N__1961\,
            I => \value_cntZ0Z_23\
        );

    \I__383\ : IoInMux
    port map (
            O => \N__1956\,
            I => \N__1953\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__1953\,
            I => \N__1950\
        );

    \I__381\ : Span4Mux_s2_h
    port map (
            O => \N__1950\,
            I => \N__1947\
        );

    \I__380\ : Span4Mux_h
    port map (
            O => \N__1947\,
            I => \N__1942\
        );

    \I__379\ : InMux
    port map (
            O => \N__1946\,
            I => \N__1937\
        );

    \I__378\ : InMux
    port map (
            O => \N__1945\,
            I => \N__1937\
        );

    \I__377\ : Odrv4
    port map (
            O => \N__1942\,
            I => leds_c_0
        );

    \I__376\ : LocalMux
    port map (
            O => \N__1937\,
            I => leds_c_0
        );

    \I__375\ : CascadeMux
    port map (
            O => \N__1932\,
            I => \N__1929\
        );

    \I__374\ : InMux
    port map (
            O => \N__1929\,
            I => \N__1922\
        );

    \I__373\ : InMux
    port map (
            O => \N__1928\,
            I => \N__1922\
        );

    \I__372\ : InMux
    port map (
            O => \N__1927\,
            I => \N__1919\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__1922\,
            I => \register10Z0Z_0\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__1919\,
            I => \register10Z0Z_0\
        );

    \I__369\ : IoInMux
    port map (
            O => \N__1914\,
            I => \N__1911\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__1911\,
            I => \N__1908\
        );

    \I__367\ : Span12Mux_s6_h
    port map (
            O => \N__1908\,
            I => \N__1903\
        );

    \I__366\ : InMux
    port map (
            O => \N__1907\,
            I => \N__1900\
        );

    \I__365\ : InMux
    port map (
            O => \N__1906\,
            I => \N__1897\
        );

    \I__364\ : Odrv12
    port map (
            O => \N__1903\,
            I => leds_c_1
        );

    \I__363\ : LocalMux
    port map (
            O => \N__1900\,
            I => leds_c_1
        );

    \I__362\ : LocalMux
    port map (
            O => \N__1897\,
            I => leds_c_1
        );

    \I__361\ : IoInMux
    port map (
            O => \N__1890\,
            I => \N__1887\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__1887\,
            I => \N__1884\
        );

    \I__359\ : Span4Mux_s2_h
    port map (
            O => \N__1884\,
            I => \N__1881\
        );

    \I__358\ : Span4Mux_h
    port map (
            O => \N__1881\,
            I => \N__1876\
        );

    \I__357\ : InMux
    port map (
            O => \N__1880\,
            I => \N__1873\
        );

    \I__356\ : InMux
    port map (
            O => \N__1879\,
            I => \N__1870\
        );

    \I__355\ : Odrv4
    port map (
            O => \N__1876\,
            I => leds_c_2
        );

    \I__354\ : LocalMux
    port map (
            O => \N__1873\,
            I => leds_c_2
        );

    \I__353\ : LocalMux
    port map (
            O => \N__1870\,
            I => leds_c_2
        );

    \I__352\ : CascadeMux
    port map (
            O => \N__1863\,
            I => \N__1858\
        );

    \I__351\ : InMux
    port map (
            O => \N__1862\,
            I => \N__1855\
        );

    \I__350\ : InMux
    port map (
            O => \N__1861\,
            I => \N__1852\
        );

    \I__349\ : InMux
    port map (
            O => \N__1858\,
            I => \N__1849\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__1855\,
            I => \value_cntZ0Z_13\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__1852\,
            I => \value_cntZ0Z_13\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__1849\,
            I => \value_cntZ0Z_13\
        );

    \I__345\ : InMux
    port map (
            O => \N__1842\,
            I => \N__1839\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__1839\,
            I => \value_cnt_cry_12_THRU_CO\
        );

    \I__343\ : InMux
    port map (
            O => \N__1836\,
            I => value_cnt_cry_12
        );

    \I__342\ : CascadeMux
    port map (
            O => \N__1833\,
            I => \N__1828\
        );

    \I__341\ : CascadeMux
    port map (
            O => \N__1832\,
            I => \N__1825\
        );

    \I__340\ : InMux
    port map (
            O => \N__1831\,
            I => \N__1822\
        );

    \I__339\ : InMux
    port map (
            O => \N__1828\,
            I => \N__1819\
        );

    \I__338\ : InMux
    port map (
            O => \N__1825\,
            I => \N__1816\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__1822\,
            I => \value_cntZ0Z_14\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__1819\,
            I => \value_cntZ0Z_14\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__1816\,
            I => \value_cntZ0Z_14\
        );

    \I__334\ : InMux
    port map (
            O => \N__1809\,
            I => \N__1806\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__1806\,
            I => \value_cnt_cry_13_THRU_CO\
        );

    \I__332\ : InMux
    port map (
            O => \N__1803\,
            I => value_cnt_cry_13
        );

    \I__331\ : CascadeMux
    port map (
            O => \N__1800\,
            I => \N__1795\
        );

    \I__330\ : InMux
    port map (
            O => \N__1799\,
            I => \N__1792\
        );

    \I__329\ : InMux
    port map (
            O => \N__1798\,
            I => \N__1789\
        );

    \I__328\ : InMux
    port map (
            O => \N__1795\,
            I => \N__1786\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__1792\,
            I => \value_cntZ0Z_15\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__1789\,
            I => \value_cntZ0Z_15\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__1786\,
            I => \value_cntZ0Z_15\
        );

    \I__324\ : InMux
    port map (
            O => \N__1779\,
            I => \N__1776\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__1776\,
            I => \value_cnt_cry_14_THRU_CO\
        );

    \I__322\ : InMux
    port map (
            O => \N__1773\,
            I => value_cnt_cry_14
        );

    \I__321\ : CascadeMux
    port map (
            O => \N__1770\,
            I => \N__1765\
        );

    \I__320\ : InMux
    port map (
            O => \N__1769\,
            I => \N__1762\
        );

    \I__319\ : InMux
    port map (
            O => \N__1768\,
            I => \N__1759\
        );

    \I__318\ : InMux
    port map (
            O => \N__1765\,
            I => \N__1756\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__1762\,
            I => \value_cntZ0Z_16\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__1759\,
            I => \value_cntZ0Z_16\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__1756\,
            I => \value_cntZ0Z_16\
        );

    \I__314\ : InMux
    port map (
            O => \N__1749\,
            I => \N__1746\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__1746\,
            I => \value_cnt_cry_15_THRU_CO\
        );

    \I__312\ : InMux
    port map (
            O => \N__1743\,
            I => \bfn_6_7_0_\
        );

    \I__311\ : CascadeMux
    port map (
            O => \N__1740\,
            I => \N__1736\
        );

    \I__310\ : InMux
    port map (
            O => \N__1739\,
            I => \N__1732\
        );

    \I__309\ : InMux
    port map (
            O => \N__1736\,
            I => \N__1729\
        );

    \I__308\ : InMux
    port map (
            O => \N__1735\,
            I => \N__1726\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__1732\,
            I => \value_cntZ0Z_17\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__1729\,
            I => \value_cntZ0Z_17\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__1726\,
            I => \value_cntZ0Z_17\
        );

    \I__304\ : InMux
    port map (
            O => \N__1719\,
            I => \N__1716\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__1716\,
            I => \value_cnt_cry_16_THRU_CO\
        );

    \I__302\ : InMux
    port map (
            O => \N__1713\,
            I => value_cnt_cry_16
        );

    \I__301\ : CascadeMux
    port map (
            O => \N__1710\,
            I => \N__1705\
        );

    \I__300\ : CascadeMux
    port map (
            O => \N__1709\,
            I => \N__1702\
        );

    \I__299\ : InMux
    port map (
            O => \N__1708\,
            I => \N__1699\
        );

    \I__298\ : InMux
    port map (
            O => \N__1705\,
            I => \N__1696\
        );

    \I__297\ : InMux
    port map (
            O => \N__1702\,
            I => \N__1693\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__1699\,
            I => \value_cntZ0Z_18\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__1696\,
            I => \value_cntZ0Z_18\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__1693\,
            I => \value_cntZ0Z_18\
        );

    \I__293\ : InMux
    port map (
            O => \N__1686\,
            I => \N__1683\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__1683\,
            I => \value_cnt_cry_17_THRU_CO\
        );

    \I__291\ : InMux
    port map (
            O => \N__1680\,
            I => value_cnt_cry_17
        );

    \I__290\ : CascadeMux
    port map (
            O => \N__1677\,
            I => \N__1673\
        );

    \I__289\ : InMux
    port map (
            O => \N__1676\,
            I => \N__1669\
        );

    \I__288\ : InMux
    port map (
            O => \N__1673\,
            I => \N__1666\
        );

    \I__287\ : InMux
    port map (
            O => \N__1672\,
            I => \N__1663\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__1669\,
            I => \value_cntZ0Z_19\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__1666\,
            I => \value_cntZ0Z_19\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__1663\,
            I => \value_cntZ0Z_19\
        );

    \I__283\ : InMux
    port map (
            O => \N__1656\,
            I => \N__1653\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__1653\,
            I => \value_cnt_cry_18_THRU_CO\
        );

    \I__281\ : InMux
    port map (
            O => \N__1650\,
            I => value_cnt_cry_18
        );

    \I__280\ : CascadeMux
    port map (
            O => \N__1647\,
            I => \N__1642\
        );

    \I__279\ : InMux
    port map (
            O => \N__1646\,
            I => \N__1639\
        );

    \I__278\ : InMux
    port map (
            O => \N__1645\,
            I => \N__1636\
        );

    \I__277\ : InMux
    port map (
            O => \N__1642\,
            I => \N__1633\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__1639\,
            I => \value_cntZ0Z_20\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__1636\,
            I => \value_cntZ0Z_20\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__1633\,
            I => \value_cntZ0Z_20\
        );

    \I__273\ : InMux
    port map (
            O => \N__1626\,
            I => \N__1623\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__1623\,
            I => \value_cnt_cry_19_THRU_CO\
        );

    \I__271\ : InMux
    port map (
            O => \N__1620\,
            I => value_cnt_cry_19
        );

    \I__270\ : CascadeMux
    port map (
            O => \N__1617\,
            I => \N__1612\
        );

    \I__269\ : InMux
    port map (
            O => \N__1616\,
            I => \N__1609\
        );

    \I__268\ : InMux
    port map (
            O => \N__1615\,
            I => \N__1606\
        );

    \I__267\ : InMux
    port map (
            O => \N__1612\,
            I => \N__1603\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__1609\,
            I => \value_cntZ0Z_5\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__1606\,
            I => \value_cntZ0Z_5\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__1603\,
            I => \value_cntZ0Z_5\
        );

    \I__263\ : InMux
    port map (
            O => \N__1596\,
            I => \N__1593\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__1593\,
            I => \value_cnt_cry_4_THRU_CO\
        );

    \I__261\ : InMux
    port map (
            O => \N__1590\,
            I => value_cnt_cry_4
        );

    \I__260\ : CascadeMux
    port map (
            O => \N__1587\,
            I => \N__1582\
        );

    \I__259\ : CascadeMux
    port map (
            O => \N__1586\,
            I => \N__1579\
        );

    \I__258\ : InMux
    port map (
            O => \N__1585\,
            I => \N__1576\
        );

    \I__257\ : InMux
    port map (
            O => \N__1582\,
            I => \N__1573\
        );

    \I__256\ : InMux
    port map (
            O => \N__1579\,
            I => \N__1570\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__1576\,
            I => \value_cntZ0Z_6\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__1573\,
            I => \value_cntZ0Z_6\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__1570\,
            I => \value_cntZ0Z_6\
        );

    \I__252\ : InMux
    port map (
            O => \N__1563\,
            I => \N__1560\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__1560\,
            I => \value_cnt_cry_5_THRU_CO\
        );

    \I__250\ : InMux
    port map (
            O => \N__1557\,
            I => value_cnt_cry_5
        );

    \I__249\ : CascadeMux
    port map (
            O => \N__1554\,
            I => \N__1549\
        );

    \I__248\ : InMux
    port map (
            O => \N__1553\,
            I => \N__1546\
        );

    \I__247\ : InMux
    port map (
            O => \N__1552\,
            I => \N__1543\
        );

    \I__246\ : InMux
    port map (
            O => \N__1549\,
            I => \N__1540\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__1546\,
            I => \value_cntZ0Z_7\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__1543\,
            I => \value_cntZ0Z_7\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__1540\,
            I => \value_cntZ0Z_7\
        );

    \I__242\ : InMux
    port map (
            O => \N__1533\,
            I => \N__1530\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__1530\,
            I => \value_cnt_cry_6_THRU_CO\
        );

    \I__240\ : InMux
    port map (
            O => \N__1527\,
            I => value_cnt_cry_6
        );

    \I__239\ : CascadeMux
    port map (
            O => \N__1524\,
            I => \N__1519\
        );

    \I__238\ : InMux
    port map (
            O => \N__1523\,
            I => \N__1516\
        );

    \I__237\ : InMux
    port map (
            O => \N__1522\,
            I => \N__1513\
        );

    \I__236\ : InMux
    port map (
            O => \N__1519\,
            I => \N__1510\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__1516\,
            I => \value_cntZ0Z_8\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__1513\,
            I => \value_cntZ0Z_8\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__1510\,
            I => \value_cntZ0Z_8\
        );

    \I__232\ : InMux
    port map (
            O => \N__1503\,
            I => \N__1500\
        );

    \I__231\ : LocalMux
    port map (
            O => \N__1500\,
            I => \value_cnt_cry_7_THRU_CO\
        );

    \I__230\ : InMux
    port map (
            O => \N__1497\,
            I => \bfn_6_6_0_\
        );

    \I__229\ : InMux
    port map (
            O => \N__1494\,
            I => value_cnt_cry_8
        );

    \I__228\ : CascadeMux
    port map (
            O => \N__1491\,
            I => \N__1486\
        );

    \I__227\ : CascadeMux
    port map (
            O => \N__1490\,
            I => \N__1483\
        );

    \I__226\ : InMux
    port map (
            O => \N__1489\,
            I => \N__1480\
        );

    \I__225\ : InMux
    port map (
            O => \N__1486\,
            I => \N__1477\
        );

    \I__224\ : InMux
    port map (
            O => \N__1483\,
            I => \N__1474\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__1480\,
            I => \value_cntZ0Z_10\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__1477\,
            I => \value_cntZ0Z_10\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__1474\,
            I => \value_cntZ0Z_10\
        );

    \I__220\ : InMux
    port map (
            O => \N__1467\,
            I => \N__1464\
        );

    \I__219\ : LocalMux
    port map (
            O => \N__1464\,
            I => \value_cnt_cry_9_THRU_CO\
        );

    \I__218\ : InMux
    port map (
            O => \N__1461\,
            I => value_cnt_cry_9
        );

    \I__217\ : InMux
    port map (
            O => \N__1458\,
            I => value_cnt_cry_10
        );

    \I__216\ : CascadeMux
    port map (
            O => \N__1455\,
            I => \N__1450\
        );

    \I__215\ : InMux
    port map (
            O => \N__1454\,
            I => \N__1447\
        );

    \I__214\ : InMux
    port map (
            O => \N__1453\,
            I => \N__1444\
        );

    \I__213\ : InMux
    port map (
            O => \N__1450\,
            I => \N__1441\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__1447\,
            I => \value_cntZ0Z_12\
        );

    \I__211\ : LocalMux
    port map (
            O => \N__1444\,
            I => \value_cntZ0Z_12\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__1441\,
            I => \value_cntZ0Z_12\
        );

    \I__209\ : InMux
    port map (
            O => \N__1434\,
            I => \N__1431\
        );

    \I__208\ : LocalMux
    port map (
            O => \N__1431\,
            I => \value_cnt_cry_11_THRU_CO\
        );

    \I__207\ : InMux
    port map (
            O => \N__1428\,
            I => value_cnt_cry_11
        );

    \I__206\ : InMux
    port map (
            O => \N__1425\,
            I => \N__1419\
        );

    \I__205\ : InMux
    port map (
            O => \N__1424\,
            I => \N__1419\
        );

    \I__204\ : LocalMux
    port map (
            O => \N__1419\,
            I => \UC.epZ0Z_0\
        );

    \I__203\ : InMux
    port map (
            O => \N__1416\,
            I => \N__1413\
        );

    \I__202\ : LocalMux
    port map (
            O => \N__1413\,
            I => \UC.epZ0Z_8\
        );

    \I__201\ : InMux
    port map (
            O => \N__1410\,
            I => \N__1404\
        );

    \I__200\ : InMux
    port map (
            O => \N__1409\,
            I => \N__1404\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__1404\,
            I => \UC.epZ0Z_1\
        );

    \I__198\ : InMux
    port map (
            O => \N__1401\,
            I => \N__1396\
        );

    \I__197\ : InMux
    port map (
            O => \N__1400\,
            I => \N__1393\
        );

    \I__196\ : InMux
    port map (
            O => \N__1399\,
            I => \N__1390\
        );

    \I__195\ : LocalMux
    port map (
            O => \N__1396\,
            I => \UC.epZ0Z_7\
        );

    \I__194\ : LocalMux
    port map (
            O => \N__1393\,
            I => \UC.epZ0Z_7\
        );

    \I__193\ : LocalMux
    port map (
            O => \N__1390\,
            I => \UC.epZ0Z_7\
        );

    \I__192\ : InMux
    port map (
            O => \N__1383\,
            I => \N__1378\
        );

    \I__191\ : InMux
    port map (
            O => \N__1382\,
            I => \N__1375\
        );

    \I__190\ : InMux
    port map (
            O => \N__1381\,
            I => \N__1372\
        );

    \I__189\ : LocalMux
    port map (
            O => \N__1378\,
            I => \value_cntZ0Z_0\
        );

    \I__188\ : LocalMux
    port map (
            O => \N__1375\,
            I => \value_cntZ0Z_0\
        );

    \I__187\ : LocalMux
    port map (
            O => \N__1372\,
            I => \value_cntZ0Z_0\
        );

    \I__186\ : CascadeMux
    port map (
            O => \N__1365\,
            I => \N__1360\
        );

    \I__185\ : InMux
    port map (
            O => \N__1364\,
            I => \N__1357\
        );

    \I__184\ : InMux
    port map (
            O => \N__1363\,
            I => \N__1354\
        );

    \I__183\ : InMux
    port map (
            O => \N__1360\,
            I => \N__1351\
        );

    \I__182\ : LocalMux
    port map (
            O => \N__1357\,
            I => \value_cntZ0Z_1\
        );

    \I__181\ : LocalMux
    port map (
            O => \N__1354\,
            I => \value_cntZ0Z_1\
        );

    \I__180\ : LocalMux
    port map (
            O => \N__1351\,
            I => \value_cntZ0Z_1\
        );

    \I__179\ : InMux
    port map (
            O => \N__1344\,
            I => \N__1341\
        );

    \I__178\ : LocalMux
    port map (
            O => \N__1341\,
            I => \value_cnt_cry_0_THRU_CO\
        );

    \I__177\ : InMux
    port map (
            O => \N__1338\,
            I => value_cnt_cry_0
        );

    \I__176\ : CascadeMux
    port map (
            O => \N__1335\,
            I => \N__1330\
        );

    \I__175\ : CascadeMux
    port map (
            O => \N__1334\,
            I => \N__1327\
        );

    \I__174\ : InMux
    port map (
            O => \N__1333\,
            I => \N__1324\
        );

    \I__173\ : InMux
    port map (
            O => \N__1330\,
            I => \N__1321\
        );

    \I__172\ : InMux
    port map (
            O => \N__1327\,
            I => \N__1318\
        );

    \I__171\ : LocalMux
    port map (
            O => \N__1324\,
            I => \value_cntZ0Z_2\
        );

    \I__170\ : LocalMux
    port map (
            O => \N__1321\,
            I => \value_cntZ0Z_2\
        );

    \I__169\ : LocalMux
    port map (
            O => \N__1318\,
            I => \value_cntZ0Z_2\
        );

    \I__168\ : InMux
    port map (
            O => \N__1311\,
            I => \N__1308\
        );

    \I__167\ : LocalMux
    port map (
            O => \N__1308\,
            I => \value_cnt_cry_1_THRU_CO\
        );

    \I__166\ : InMux
    port map (
            O => \N__1305\,
            I => value_cnt_cry_1
        );

    \I__165\ : CascadeMux
    port map (
            O => \N__1302\,
            I => \N__1297\
        );

    \I__164\ : InMux
    port map (
            O => \N__1301\,
            I => \N__1294\
        );

    \I__163\ : InMux
    port map (
            O => \N__1300\,
            I => \N__1291\
        );

    \I__162\ : InMux
    port map (
            O => \N__1297\,
            I => \N__1288\
        );

    \I__161\ : LocalMux
    port map (
            O => \N__1294\,
            I => \value_cntZ0Z_3\
        );

    \I__160\ : LocalMux
    port map (
            O => \N__1291\,
            I => \value_cntZ0Z_3\
        );

    \I__159\ : LocalMux
    port map (
            O => \N__1288\,
            I => \value_cntZ0Z_3\
        );

    \I__158\ : InMux
    port map (
            O => \N__1281\,
            I => \N__1278\
        );

    \I__157\ : LocalMux
    port map (
            O => \N__1278\,
            I => \value_cnt_cry_2_THRU_CO\
        );

    \I__156\ : InMux
    port map (
            O => \N__1275\,
            I => value_cnt_cry_2
        );

    \I__155\ : CascadeMux
    port map (
            O => \N__1272\,
            I => \N__1267\
        );

    \I__154\ : InMux
    port map (
            O => \N__1271\,
            I => \N__1264\
        );

    \I__153\ : InMux
    port map (
            O => \N__1270\,
            I => \N__1261\
        );

    \I__152\ : InMux
    port map (
            O => \N__1267\,
            I => \N__1258\
        );

    \I__151\ : LocalMux
    port map (
            O => \N__1264\,
            I => \value_cntZ0Z_4\
        );

    \I__150\ : LocalMux
    port map (
            O => \N__1261\,
            I => \value_cntZ0Z_4\
        );

    \I__149\ : LocalMux
    port map (
            O => \N__1258\,
            I => \value_cntZ0Z_4\
        );

    \I__148\ : InMux
    port map (
            O => \N__1251\,
            I => \N__1248\
        );

    \I__147\ : LocalMux
    port map (
            O => \N__1248\,
            I => \value_cnt_cry_3_THRU_CO\
        );

    \I__146\ : InMux
    port map (
            O => \N__1245\,
            I => value_cnt_cry_3
        );

    \I__145\ : InMux
    port map (
            O => \N__1242\,
            I => \N__1237\
        );

    \I__144\ : InMux
    port map (
            O => \N__1241\,
            I => \N__1234\
        );

    \I__143\ : InMux
    port map (
            O => \N__1240\,
            I => \N__1231\
        );

    \I__142\ : LocalMux
    port map (
            O => \N__1237\,
            I => \UC.epZ0Z_4\
        );

    \I__141\ : LocalMux
    port map (
            O => \N__1234\,
            I => \UC.epZ0Z_4\
        );

    \I__140\ : LocalMux
    port map (
            O => \N__1231\,
            I => \UC.epZ0Z_4\
        );

    \I__139\ : InMux
    port map (
            O => \N__1224\,
            I => \N__1220\
        );

    \I__138\ : InMux
    port map (
            O => \N__1223\,
            I => \N__1217\
        );

    \I__137\ : LocalMux
    port map (
            O => \N__1220\,
            I => \UC.sr_reg\
        );

    \I__136\ : LocalMux
    port map (
            O => \N__1217\,
            I => \UC.sr_reg\
        );

    \I__135\ : CascadeMux
    port map (
            O => \N__1212\,
            I => \N__1207\
        );

    \I__134\ : CascadeMux
    port map (
            O => \N__1211\,
            I => \N__1204\
        );

    \I__133\ : InMux
    port map (
            O => \N__1210\,
            I => \N__1194\
        );

    \I__132\ : InMux
    port map (
            O => \N__1207\,
            I => \N__1194\
        );

    \I__131\ : InMux
    port map (
            O => \N__1204\,
            I => \N__1194\
        );

    \I__130\ : InMux
    port map (
            O => \N__1203\,
            I => \N__1194\
        );

    \I__129\ : LocalMux
    port map (
            O => \N__1194\,
            I => op_eq_un4_fin_cnt_20
        );

    \I__128\ : CascadeMux
    port map (
            O => \N__1191\,
            I => \N__1186\
        );

    \I__127\ : InMux
    port map (
            O => \N__1190\,
            I => \N__1180\
        );

    \I__126\ : InMux
    port map (
            O => \N__1189\,
            I => \N__1180\
        );

    \I__125\ : InMux
    port map (
            O => \N__1186\,
            I => \N__1175\
        );

    \I__124\ : InMux
    port map (
            O => \N__1185\,
            I => \N__1175\
        );

    \I__123\ : LocalMux
    port map (
            O => \N__1180\,
            I => op_eq_un4_fin_cnt_21
        );

    \I__122\ : LocalMux
    port map (
            O => \N__1175\,
            I => op_eq_un4_fin_cnt_21
        );

    \I__121\ : InMux
    port map (
            O => \N__1170\,
            I => \N__1163\
        );

    \I__120\ : InMux
    port map (
            O => \N__1169\,
            I => \N__1163\
        );

    \I__119\ : InMux
    port map (
            O => \N__1168\,
            I => \N__1160\
        );

    \I__118\ : LocalMux
    port map (
            O => \N__1163\,
            I => \UC.epZ0Z_3\
        );

    \I__117\ : LocalMux
    port map (
            O => \N__1160\,
            I => \UC.epZ0Z_3\
        );

    \I__116\ : CascadeMux
    port map (
            O => \N__1155\,
            I => \N__1150\
        );

    \I__115\ : InMux
    port map (
            O => \N__1154\,
            I => \N__1145\
        );

    \I__114\ : InMux
    port map (
            O => \N__1153\,
            I => \N__1145\
        );

    \I__113\ : InMux
    port map (
            O => \N__1150\,
            I => \N__1142\
        );

    \I__112\ : LocalMux
    port map (
            O => \N__1145\,
            I => \UC.epZ0Z_6\
        );

    \I__111\ : LocalMux
    port map (
            O => \N__1142\,
            I => \UC.epZ0Z_6\
        );

    \I__110\ : IoInMux
    port map (
            O => \N__1137\,
            I => \N__1134\
        );

    \I__109\ : LocalMux
    port map (
            O => \N__1134\,
            I => \N__1131\
        );

    \I__108\ : Span4Mux_s0_h
    port map (
            O => \N__1131\,
            I => \N__1128\
        );

    \I__107\ : Odrv4
    port map (
            O => \N__1128\,
            I => \UC.value_cnte_0_i\
        );

    \I__106\ : CascadeMux
    port map (
            O => \N__1125\,
            I => \op_eq_un4_fin_cnt_20_3_cascade_\
        );

    \I__105\ : InMux
    port map (
            O => \N__1122\,
            I => \N__1119\
        );

    \I__104\ : LocalMux
    port map (
            O => \N__1119\,
            I => op_eq_un4_fin_cnt_20_4
        );

    \I__103\ : InMux
    port map (
            O => \N__1116\,
            I => \N__1113\
        );

    \I__102\ : LocalMux
    port map (
            O => \N__1113\,
            I => op_eq_un4_fin_cnt_21_9
        );

    \I__101\ : InMux
    port map (
            O => \N__1110\,
            I => \N__1107\
        );

    \I__100\ : LocalMux
    port map (
            O => \N__1107\,
            I => op_eq_un4_fin_cnt_21_11
        );

    \I__99\ : CascadeMux
    port map (
            O => \N__1104\,
            I => \N__1101\
        );

    \I__98\ : InMux
    port map (
            O => \N__1101\,
            I => \N__1098\
        );

    \I__97\ : LocalMux
    port map (
            O => \N__1098\,
            I => op_eq_un4_fin_cnt_21_10
        );

    \I__96\ : InMux
    port map (
            O => \N__1095\,
            I => \N__1092\
        );

    \I__95\ : LocalMux
    port map (
            O => \N__1092\,
            I => op_eq_un4_fin_cnt_21_8
        );

    \IN_MUX_bfv_6_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_5_0_\
        );

    \IN_MUX_bfv_6_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => value_cnt_cry_7,
            carryinitout => \bfn_6_6_0_\
        );

    \IN_MUX_bfv_6_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => value_cnt_cry_15,
            carryinitout => \bfn_6_7_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \UC.ep_RNI0P1C_0_3\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__1137\,
            GLOBALBUFFEROUTPUT => value_cnte_0_i_g
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \value_cnt_RNIOUPL1_8_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2142\,
            in1 => \N__1522\,
            in2 => \N__1491\,
            in3 => \N__2277\,
            lcout => op_eq_un4_fin_cnt_21_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_RNIMPFN1_12_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1861\,
            in1 => \N__1453\,
            in2 => \N__1833\,
            in3 => \N__1798\,
            lcout => op_eq_un4_fin_cnt_21_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_RNIQ34K1_4_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1615\,
            in1 => \N__1270\,
            in2 => \N__1587\,
            in3 => \N__1552\,
            lcout => op_eq_un4_fin_cnt_21_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_RNIAJ3K1_0_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1363\,
            in1 => \N__1382\,
            in2 => \N__1335\,
            in3 => \N__1300\,
            lcout => op_eq_un4_fin_cnt_21_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_RNI6AGN1_16_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1735\,
            in1 => \N__1768\,
            in2 => \N__1709\,
            in3 => \N__1672\,
            lcout => op_eq_un4_fin_cnt_20_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_RNINQPR_20_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1645\,
            in2 => \_gnd_net_\,
            in3 => \N__2026\,
            lcout => OPEN,
            ltout => \op_eq_un4_fin_cnt_20_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_RNIO34F3_23_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__1971\,
            in1 => \N__1999\,
            in2 => \N__1125\,
            in3 => \N__1122\,
            lcout => op_eq_un4_fin_cnt_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_RNIIFHL6_0_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1116\,
            in1 => \N__1110\,
            in2 => \N__1104\,
            in3 => \N__1095\,
            lcout => op_eq_un4_fin_cnt_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \UC.ep_3_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101001100"
        )
    port map (
            in0 => \N__1189\,
            in1 => \N__1169\,
            in2 => \N__1212\,
            in3 => \N__1242\,
            lcout => \UC.epZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2110\,
            ce => 'H',
            sr => \N__2063\
        );

    \UC.ep_6_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111011101110"
        )
    port map (
            in0 => \N__1154\,
            in1 => \N__1401\,
            in2 => \N__1191\,
            in3 => \N__1210\,
            lcout => \UC.epZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2110\,
            ce => 'H',
            sr => \N__2063\
        );

    \UC.ep_2_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__1170\,
            in1 => \N__1190\,
            in2 => \_gnd_net_\,
            in3 => \N__1203\,
            lcout => \UC.sr_reg\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2110\,
            ce => 'H',
            sr => \N__2063\
        );

    \UC.ep_5_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1153\,
            in2 => \N__1211\,
            in3 => \N__1185\,
            lcout => sl_reg,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2110\,
            ce => 'H',
            sr => \N__2063\
        );

    \UC.ep_RNI0P1C_3_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__1168\,
            in1 => \N__1240\,
            in2 => \N__1155\,
            in3 => \N__1399\,
            lcout => \UC.value_cnte_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_1_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__1364\,
            in1 => \N__2240\,
            in2 => \_gnd_net_\,
            in3 => \N__1344\,
            lcout => \value_cntZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2117\,
            ce => \N__2084\,
            sr => \N__2056\
        );

    \value_cnt_6_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__2245\,
            in1 => \N__1585\,
            in2 => \_gnd_net_\,
            in3 => \N__1563\,
            lcout => \value_cntZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2117\,
            ce => \N__2084\,
            sr => \N__2056\
        );

    \value_cnt_7_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__1553\,
            in1 => \N__2246\,
            in2 => \_gnd_net_\,
            in3 => \N__1533\,
            lcout => \value_cntZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2117\,
            ce => \N__2084\,
            sr => \N__2056\
        );

    \value_cnt_4_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__2243\,
            in1 => \N__1271\,
            in2 => \_gnd_net_\,
            in3 => \N__1251\,
            lcout => \value_cntZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2117\,
            ce => \N__2084\,
            sr => \N__2056\
        );

    \value_cnt_3_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__1301\,
            in1 => \N__2242\,
            in2 => \_gnd_net_\,
            in3 => \N__1281\,
            lcout => \value_cntZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2117\,
            ce => \N__2084\,
            sr => \N__2056\
        );

    \value_cnt_2_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__2241\,
            in1 => \N__1333\,
            in2 => \_gnd_net_\,
            in3 => \N__1311\,
            lcout => \value_cntZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2117\,
            ce => \N__2084\,
            sr => \N__2056\
        );

    \value_cnt_5_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__1616\,
            in1 => \N__2244\,
            in2 => \_gnd_net_\,
            in3 => \N__1596\,
            lcout => \value_cntZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2117\,
            ce => \N__2084\,
            sr => \N__2056\
        );

    \value_cnt_14_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__2237\,
            in1 => \N__1831\,
            in2 => \_gnd_net_\,
            in3 => \N__1809\,
            lcout => \value_cntZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2114\,
            ce => \N__2082\,
            sr => \N__2058\
        );

    \value_cnt_10_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__2234\,
            in1 => \N__1489\,
            in2 => \_gnd_net_\,
            in3 => \N__1467\,
            lcout => \value_cntZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2114\,
            ce => \N__2082\,
            sr => \N__2058\
        );

    \value_cnt_0_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2233\,
            in2 => \_gnd_net_\,
            in3 => \N__1383\,
            lcout => \value_cntZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2114\,
            ce => \N__2082\,
            sr => \N__2058\
        );

    \value_cnt_8_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__2239\,
            in1 => \N__1523\,
            in2 => \_gnd_net_\,
            in3 => \N__1503\,
            lcout => \value_cntZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2114\,
            ce => \N__2082\,
            sr => \N__2058\
        );

    \value_cnt_13_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__1862\,
            in1 => \N__2236\,
            in2 => \_gnd_net_\,
            in3 => \N__1842\,
            lcout => \value_cntZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2114\,
            ce => \N__2082\,
            sr => \N__2058\
        );

    \value_cnt_12_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__2235\,
            in1 => \N__1454\,
            in2 => \_gnd_net_\,
            in3 => \N__1434\,
            lcout => \value_cntZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2114\,
            ce => \N__2082\,
            sr => \N__2058\
        );

    \value_cnt_15_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__1799\,
            in1 => \N__2238\,
            in2 => \_gnd_net_\,
            in3 => \N__1779\,
            lcout => \value_cntZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2114\,
            ce => \N__2082\,
            sr => \N__2058\
        );

    \value_cnt_18_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__2193\,
            in1 => \N__1708\,
            in2 => \_gnd_net_\,
            in3 => \N__1686\,
            lcout => \value_cntZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2112\,
            ce => \N__2081\,
            sr => \N__2061\
        );

    \value_cnt_22_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__2001\,
            in1 => \N__2196\,
            in2 => \_gnd_net_\,
            in3 => \N__1983\,
            lcout => \value_cntZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2112\,
            ce => \N__2081\,
            sr => \N__2061\
        );

    \value_cnt_19_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__2194\,
            in1 => \N__1676\,
            in2 => \_gnd_net_\,
            in3 => \N__1656\,
            lcout => \value_cntZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2112\,
            ce => \N__2081\,
            sr => \N__2061\
        );

    \value_cnt_20_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__2195\,
            in1 => \N__1646\,
            in2 => \_gnd_net_\,
            in3 => \N__1626\,
            lcout => \value_cntZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2112\,
            ce => \N__2081\,
            sr => \N__2061\
        );

    \value_cnt_17_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__2197\,
            in1 => \N__1739\,
            in2 => \_gnd_net_\,
            in3 => \N__1719\,
            lcout => \value_cntZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2112\,
            ce => \N__2081\,
            sr => \N__2061\
        );

    \value_cnt_16_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__2192\,
            in1 => \N__1769\,
            in2 => \_gnd_net_\,
            in3 => \N__1749\,
            lcout => \value_cntZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2112\,
            ce => \N__2081\,
            sr => \N__2061\
        );

    \value_cnt_21_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__2198\,
            in1 => \N__2030\,
            in2 => \_gnd_net_\,
            in3 => \N__2010\,
            lcout => \value_cntZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2112\,
            ce => \N__2081\,
            sr => \N__2061\
        );

    \UC.ep_RNIHT06_4_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1400\,
            in2 => \_gnd_net_\,
            in3 => \N__1241\,
            lcout => \UC_un1_ld_cnt_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \UC.ep_RNIDP06_2_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1223\,
            in2 => \_gnd_net_\,
            in3 => \N__2490\,
            lcout => un1_sr_reg_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \UC.ep_4_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__2469\,
            in1 => \N__1424\,
            in2 => \N__1932\,
            in3 => \N__1410\,
            lcout => \UC.epZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2113\,
            ce => 'H',
            sr => \N__2064\
        );

    \UC.ep_0_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1224\,
            lcout => \UC.epZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2113\,
            ce => 'H',
            sr => \N__2064\
        );

    \UC.ep_8_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__1425\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1928\,
            lcout => \UC.epZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2113\,
            ce => 'H',
            sr => \N__2064\
        );

    \UC.ep_1_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2501\,
            lcout => \UC.epZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2113\,
            ce => 'H',
            sr => \N__2064\
        );

    \UC.ep_7_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__2468\,
            in1 => \N__1416\,
            in2 => \_gnd_net_\,
            in3 => \N__1409\,
            lcout => \UC.epZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2113\,
            ce => 'H',
            sr => \N__2064\
        );

    \value_cnt_cry_c_0_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1381\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_5_0_\,
            carryout => value_cnt_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_0_THRU_LUT4_0_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2336\,
            in2 => \N__1365\,
            in3 => \N__1338\,
            lcout => \value_cnt_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_0,
            carryout => value_cnt_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_1_THRU_LUT4_0_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2340\,
            in2 => \N__1334\,
            in3 => \N__1305\,
            lcout => \value_cnt_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_1,
            carryout => value_cnt_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_2_THRU_LUT4_0_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2337\,
            in2 => \N__1302\,
            in3 => \N__1275\,
            lcout => \value_cnt_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_2,
            carryout => value_cnt_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_3_THRU_LUT4_0_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2341\,
            in2 => \N__1272\,
            in3 => \N__1245\,
            lcout => \value_cnt_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_3,
            carryout => value_cnt_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_4_THRU_LUT4_0_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2338\,
            in2 => \N__1617\,
            in3 => \N__1590\,
            lcout => \value_cnt_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_4,
            carryout => value_cnt_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_5_THRU_LUT4_0_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2342\,
            in2 => \N__1586\,
            in3 => \N__1557\,
            lcout => \value_cnt_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_5,
            carryout => value_cnt_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_6_THRU_LUT4_0_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2339\,
            in2 => \N__1554\,
            in3 => \N__1527\,
            lcout => \value_cnt_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_6,
            carryout => value_cnt_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_7_THRU_LUT4_0_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2349\,
            in2 => \N__1524\,
            in3 => \N__1497\,
            lcout => \value_cnt_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_6_6_0_\,
            carryout => value_cnt_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_8_THRU_LUT4_0_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2346\,
            in2 => \N__2141\,
            in3 => \N__1494\,
            lcout => \value_cnt_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_8,
            carryout => value_cnt_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_9_THRU_LUT4_0_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2350\,
            in2 => \N__1490\,
            in3 => \N__1461\,
            lcout => \value_cnt_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_9,
            carryout => value_cnt_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_10_THRU_LUT4_0_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2343\,
            in2 => \N__2276\,
            in3 => \N__1458\,
            lcout => \value_cnt_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_10,
            carryout => value_cnt_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_11_THRU_LUT4_0_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2347\,
            in2 => \N__1455\,
            in3 => \N__1428\,
            lcout => \value_cnt_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_11,
            carryout => value_cnt_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_12_THRU_LUT4_0_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2344\,
            in2 => \N__1863\,
            in3 => \N__1836\,
            lcout => \value_cnt_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_12,
            carryout => value_cnt_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_13_THRU_LUT4_0_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2348\,
            in2 => \N__1832\,
            in3 => \N__1803\,
            lcout => \value_cnt_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_13,
            carryout => value_cnt_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_14_THRU_LUT4_0_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2345\,
            in2 => \N__1800\,
            in3 => \N__1773\,
            lcout => \value_cnt_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_14,
            carryout => value_cnt_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_15_THRU_LUT4_0_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2376\,
            in2 => \N__1770\,
            in3 => \N__1743\,
            lcout => \value_cnt_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_6_7_0_\,
            carryout => value_cnt_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_16_THRU_LUT4_0_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2370\,
            in2 => \N__1740\,
            in3 => \N__1713\,
            lcout => \value_cnt_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_16,
            carryout => value_cnt_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_17_THRU_LUT4_0_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2377\,
            in2 => \N__1710\,
            in3 => \N__1680\,
            lcout => \value_cnt_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_17,
            carryout => value_cnt_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_18_THRU_LUT4_0_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2371\,
            in2 => \N__1677\,
            in3 => \N__1650\,
            lcout => \value_cnt_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_18,
            carryout => value_cnt_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_19_THRU_LUT4_0_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2378\,
            in2 => \N__1647\,
            in3 => \N__1620\,
            lcout => \value_cnt_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_19,
            carryout => value_cnt_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_20_THRU_LUT4_0_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2372\,
            in2 => \N__2031\,
            in3 => \N__2004\,
            lcout => \value_cnt_cry_20_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_20,
            carryout => value_cnt_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_cry_21_THRU_LUT4_0_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2000\,
            in2 => \N__2379\,
            in3 => \N__1977\,
            lcout => \value_cnt_cry_21_THRU_CO\,
            ltout => OPEN,
            carryin => value_cnt_cry_21,
            carryout => value_cnt_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_23_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__1970\,
            in1 => \N__2214\,
            in2 => \_gnd_net_\,
            in3 => \N__1974\,
            lcout => \value_cntZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2115\,
            ce => \N__2083\,
            sr => \N__2057\
        );

    \register10_1_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__2503\,
            in1 => \N__1927\,
            in2 => \_gnd_net_\,
            in3 => \N__1906\,
            lcout => leds_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2111\,
            ce => \N__2396\,
            sr => \N__2060\
        );

    \register10_2_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__1946\,
            in1 => \N__1880\,
            in2 => \_gnd_net_\,
            in3 => \N__2504\,
            lcout => leds_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2111\,
            ce => \N__2396\,
            sr => \N__2060\
        );

    \register10_0_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__1945\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2502\,
            lcout => \register10Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2111\,
            ce => \N__2396\,
            sr => \N__2060\
        );

    \register10_3_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__2521\,
            in1 => \_gnd_net_\,
            in2 => \N__2594\,
            in3 => \N__1907\,
            lcout => leds_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2116\,
            ce => \N__2403\,
            sr => \N__2062\
        );

    \register10_6_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2447\,
            in1 => \N__2563\,
            in2 => \_gnd_net_\,
            in3 => \N__2524\,
            lcout => leds_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2116\,
            ce => \N__2403\,
            sr => \N__2062\
        );

    \register10_4_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__2522\,
            in1 => \_gnd_net_\,
            in2 => \N__2570\,
            in3 => \N__1879\,
            lcout => leds_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2116\,
            ce => \N__2403\,
            sr => \N__2062\
        );

    \register10_5_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2540\,
            in1 => \N__2587\,
            in2 => \_gnd_net_\,
            in3 => \N__2523\,
            lcout => leds_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2116\,
            ce => \N__2403\,
            sr => \N__2062\
        );

    \register10_7_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__2525\,
            in1 => \_gnd_net_\,
            in2 => \N__2423\,
            in3 => \N__2539\,
            lcout => leds_c_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2116\,
            ce => \N__2403\,
            sr => \N__2062\
        );

    \register10_9_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2416\,
            in2 => \_gnd_net_\,
            in3 => \N__2520\,
            lcout => \register10Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2116\,
            ce => \N__2403\,
            sr => \N__2062\
        );

    \register10_8_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__2526\,
            in1 => \N__2467\,
            in2 => \_gnd_net_\,
            in3 => \N__2446\,
            lcout => leds_c_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2116\,
            ce => \N__2403\,
            sr => \N__2062\
        );

    \CONSTANT_ONE_LUT4_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \value_cnt_11_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111010111011"
        )
    port map (
            in0 => \N__2252\,
            in1 => \N__2275\,
            in2 => \_gnd_net_\,
            in3 => \N__2283\,
            lcout => \value_cntZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2118\,
            ce => \N__2085\,
            sr => \N__2059\
        );

    \value_cnt_9_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101010101111"
        )
    port map (
            in0 => \N__2253\,
            in1 => \_gnd_net_\,
            in2 => \N__2151\,
            in3 => \N__2140\,
            lcout => \value_cntZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2118\,
            ce => \N__2085\,
            sr => \N__2059\
        );
end \INTERFACE\;
